//[UHDL]Content Start [md5:3634c664f0cae32a29033e3a1552312c]
module filter_subpredecoder_type_first (
	input  [31:0]  pred_pc      ,
	input  [8:0]   v_vld        ,
	input  [8:0]   v_ena        ,
	input  [8:0]   v_inst_type  ,
	input  [143:0] data         ,
	output [255:0] v_dec_inst   ,
	output [7:0]   v_dec_ena    ,
	output [7:0]   v_dec_last   ,
	output [255:0] v_dec_pc     ,
	output [255:0] v_dec_nxt_pc ,
	output         need_last_buf,
	output         use_last     );

	//Wire define for this module.
	wire [7:0]  v_dec_vld     ;
	reg  [31:0] v_dec_inst_0  ;
	reg  [0:0]  v_dec_ena_0   ;
	reg  [0:0]  v_dec_vld_0   ;
	reg  [32:0] v_dec_pc_add_0;
	reg  [31:0] v_dec_inst_1  ;
	reg  [0:0]  v_dec_ena_1   ;
	reg  [0:0]  v_dec_vld_1   ;
	reg  [32:0] v_dec_pc_add_1;
	reg  [31:0] v_dec_inst_2  ;
	reg  [0:0]  v_dec_ena_2   ;
	reg  [0:0]  v_dec_vld_2   ;
	reg  [32:0] v_dec_pc_add_2;
	reg  [31:0] v_dec_inst_3  ;
	reg  [0:0]  v_dec_ena_3   ;
	reg  [0:0]  v_dec_vld_3   ;
	reg  [32:0] v_dec_pc_add_3;
	reg  [31:0] v_dec_inst_4  ;
	reg  [0:0]  v_dec_ena_4   ;
	reg  [0:0]  v_dec_vld_4   ;
	reg  [32:0] v_dec_pc_add_4;
	reg  [31:0] v_dec_inst_5  ;
	reg  [0:0]  v_dec_ena_5   ;
	reg  [0:0]  v_dec_vld_5   ;
	reg  [32:0] v_dec_pc_add_5;
	reg  [31:0] v_dec_inst_6  ;
	reg  [0:0]  v_dec_ena_6   ;
	reg  [0:0]  v_dec_vld_6   ;
	reg  [32:0] v_dec_pc_add_6;
	reg  [31:0] v_dec_inst_7  ;
	reg  [0:0]  v_dec_ena_7   ;
	reg  [0:0]  v_dec_vld_7   ;
	reg  [32:0] v_dec_pc_add_7;
	reg  [0:0]  use_last_w    ;

	//Wire define for sub module.

	//Wire define for Inout.

	//Wire sub module connect to this module and inter module connect.
	assign v_dec_inst = {v_dec_inst_7, v_dec_inst_6, v_dec_inst_5, v_dec_inst_4, v_dec_inst_3, v_dec_inst_2, v_dec_inst_1, v_dec_inst_0};
	
	assign v_dec_ena = {v_dec_ena_7, v_dec_ena_6, v_dec_ena_5, v_dec_ena_4, v_dec_ena_3, v_dec_ena_2, v_dec_ena_1, v_dec_ena_0};
	
	assign v_dec_pc = {v_dec_pc_add_6[31:0], v_dec_pc_add_5[31:0], v_dec_pc_add_4[31:0], v_dec_pc_add_3[31:0], v_dec_pc_add_2[31:0], v_dec_pc_add_1[31:0], v_dec_pc_add_0[31:0], pred_pc};
	
	assign v_dec_nxt_pc = {v_dec_pc_add_7[31:0], v_dec_pc_add_6[31:0], v_dec_pc_add_5[31:0], v_dec_pc_add_4[31:0], v_dec_pc_add_3[31:0], v_dec_pc_add_2[31:0], v_dec_pc_add_1[31:0], v_dec_pc_add_0[31:0]};
	
	assign need_last_buf = ((|v_dec_vld) && (!(&v_vld)));
	
	assign use_last = use_last_w;
	
	assign v_dec_vld = {v_dec_vld_7, v_dec_vld_6, v_dec_vld_5, v_dec_vld_4, v_dec_vld_3, v_dec_vld_2, v_dec_vld_1, v_dec_vld_0};
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_inst_0 = data[31:0];
	    8'b1111110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1111101 : v_dec_inst_0 = data[31:0];
	    8'b1111100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1111011 : v_dec_inst_0 = data[31:0];
	    8'b1111010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1111001 : v_dec_inst_0 = data[31:0];
	    8'b1111000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1110111 : v_dec_inst_0 = data[31:0];
	    8'b1110110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1110101 : v_dec_inst_0 = data[31:0];
	    8'b1110100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1110011 : v_dec_inst_0 = data[31:0];
	    8'b1110010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1110001 : v_dec_inst_0 = data[31:0];
	    8'b1110000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1101111 : v_dec_inst_0 = data[31:0];
	    8'b1101110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1101101 : v_dec_inst_0 = data[31:0];
	    8'b1101100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1101011 : v_dec_inst_0 = data[31:0];
	    8'b1101010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1101001 : v_dec_inst_0 = data[31:0];
	    8'b1101000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1100111 : v_dec_inst_0 = data[31:0];
	    8'b1100110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1100101 : v_dec_inst_0 = data[31:0];
	    8'b1100100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1100011 : v_dec_inst_0 = data[31:0];
	    8'b1100010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1100001 : v_dec_inst_0 = data[31:0];
	    8'b1100000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1011111 : v_dec_inst_0 = data[31:0];
	    8'b1011110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1011101 : v_dec_inst_0 = data[31:0];
	    8'b1011100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1011011 : v_dec_inst_0 = data[31:0];
	    8'b1011010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1011001 : v_dec_inst_0 = data[31:0];
	    8'b1011000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1010111 : v_dec_inst_0 = data[31:0];
	    8'b1010110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1010101 : v_dec_inst_0 = data[31:0];
	    8'b1010100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1010011 : v_dec_inst_0 = data[31:0];
	    8'b1010010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1010001 : v_dec_inst_0 = data[31:0];
	    8'b1010000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1001111 : v_dec_inst_0 = data[31:0];
	    8'b1001110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1001101 : v_dec_inst_0 = data[31:0];
	    8'b1001100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1001011 : v_dec_inst_0 = data[31:0];
	    8'b1001010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1001001 : v_dec_inst_0 = data[31:0];
	    8'b1001000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1000111 : v_dec_inst_0 = data[31:0];
	    8'b1000110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1000101 : v_dec_inst_0 = data[31:0];
	    8'b1000100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1000011 : v_dec_inst_0 = data[31:0];
	    8'b1000010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1000001 : v_dec_inst_0 = data[31:0];
	    8'b1000000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b111111 : v_dec_inst_0 = data[31:0];
	    8'b111110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b111101 : v_dec_inst_0 = data[31:0];
	    8'b111100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b111011 : v_dec_inst_0 = data[31:0];
	    8'b111010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b111001 : v_dec_inst_0 = data[31:0];
	    8'b111000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b110111 : v_dec_inst_0 = data[31:0];
	    8'b110110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b110101 : v_dec_inst_0 = data[31:0];
	    8'b110100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b110011 : v_dec_inst_0 = data[31:0];
	    8'b110010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b110001 : v_dec_inst_0 = data[31:0];
	    8'b110000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b101111 : v_dec_inst_0 = data[31:0];
	    8'b101110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b101101 : v_dec_inst_0 = data[31:0];
	    8'b101100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b101011 : v_dec_inst_0 = data[31:0];
	    8'b101010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b101001 : v_dec_inst_0 = data[31:0];
	    8'b101000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b100111 : v_dec_inst_0 = data[31:0];
	    8'b100110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b100101 : v_dec_inst_0 = data[31:0];
	    8'b100100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b100011 : v_dec_inst_0 = data[31:0];
	    8'b100010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b100001 : v_dec_inst_0 = data[31:0];
	    8'b100000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11111 : v_dec_inst_0 = data[31:0];
	    8'b11110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11101 : v_dec_inst_0 = data[31:0];
	    8'b11100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11011 : v_dec_inst_0 = data[31:0];
	    8'b11010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11001 : v_dec_inst_0 = data[31:0];
	    8'b11000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10111 : v_dec_inst_0 = data[31:0];
	    8'b10110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10101 : v_dec_inst_0 = data[31:0];
	    8'b10100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10011 : v_dec_inst_0 = data[31:0];
	    8'b10010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10001 : v_dec_inst_0 = data[31:0];
	    8'b10000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1111 : v_dec_inst_0 = data[31:0];
	    8'b1110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1101 : v_dec_inst_0 = data[31:0];
	    8'b1100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1011 : v_dec_inst_0 = data[31:0];
	    8'b1010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1001 : v_dec_inst_0 = data[31:0];
	    8'b1000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b111 : v_dec_inst_0 = data[31:0];
	    8'b110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b101 : v_dec_inst_0 = data[31:0];
	    8'b100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11 : v_dec_inst_0 = data[31:0];
	    8'b10 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b1 : v_dec_inst_0 = data[31:0];
	    8'b0 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11111111 : v_dec_inst_0 = data[31:0];
	    8'b11111110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11111101 : v_dec_inst_0 = data[31:0];
	    8'b11111100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11111011 : v_dec_inst_0 = data[31:0];
	    8'b11111010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11111001 : v_dec_inst_0 = data[31:0];
	    8'b11111000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11110111 : v_dec_inst_0 = data[31:0];
	    8'b11110110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11110101 : v_dec_inst_0 = data[31:0];
	    8'b11110100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11110011 : v_dec_inst_0 = data[31:0];
	    8'b11110010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11110001 : v_dec_inst_0 = data[31:0];
	    8'b11110000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11101111 : v_dec_inst_0 = data[31:0];
	    8'b11101110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11101101 : v_dec_inst_0 = data[31:0];
	    8'b11101100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11101011 : v_dec_inst_0 = data[31:0];
	    8'b11101010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11101001 : v_dec_inst_0 = data[31:0];
	    8'b11101000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11100111 : v_dec_inst_0 = data[31:0];
	    8'b11100110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11100101 : v_dec_inst_0 = data[31:0];
	    8'b11100100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11100011 : v_dec_inst_0 = data[31:0];
	    8'b11100010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11100001 : v_dec_inst_0 = data[31:0];
	    8'b11100000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11011111 : v_dec_inst_0 = data[31:0];
	    8'b11011110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11011101 : v_dec_inst_0 = data[31:0];
	    8'b11011100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11011011 : v_dec_inst_0 = data[31:0];
	    8'b11011010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11011001 : v_dec_inst_0 = data[31:0];
	    8'b11011000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11010111 : v_dec_inst_0 = data[31:0];
	    8'b11010110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11010101 : v_dec_inst_0 = data[31:0];
	    8'b11010100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11010011 : v_dec_inst_0 = data[31:0];
	    8'b11010010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11010001 : v_dec_inst_0 = data[31:0];
	    8'b11010000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11001111 : v_dec_inst_0 = data[31:0];
	    8'b11001110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11001101 : v_dec_inst_0 = data[31:0];
	    8'b11001100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11001011 : v_dec_inst_0 = data[31:0];
	    8'b11001010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11001001 : v_dec_inst_0 = data[31:0];
	    8'b11001000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11000111 : v_dec_inst_0 = data[31:0];
	    8'b11000110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11000101 : v_dec_inst_0 = data[31:0];
	    8'b11000100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11000011 : v_dec_inst_0 = data[31:0];
	    8'b11000010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b11000001 : v_dec_inst_0 = data[31:0];
	    8'b11000000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10111111 : v_dec_inst_0 = data[31:0];
	    8'b10111110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10111101 : v_dec_inst_0 = data[31:0];
	    8'b10111100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10111011 : v_dec_inst_0 = data[31:0];
	    8'b10111010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10111001 : v_dec_inst_0 = data[31:0];
	    8'b10111000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10110111 : v_dec_inst_0 = data[31:0];
	    8'b10110110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10110101 : v_dec_inst_0 = data[31:0];
	    8'b10110100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10110011 : v_dec_inst_0 = data[31:0];
	    8'b10110010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10110001 : v_dec_inst_0 = data[31:0];
	    8'b10110000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10101111 : v_dec_inst_0 = data[31:0];
	    8'b10101110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10101101 : v_dec_inst_0 = data[31:0];
	    8'b10101100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10101011 : v_dec_inst_0 = data[31:0];
	    8'b10101010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10101001 : v_dec_inst_0 = data[31:0];
	    8'b10101000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10100111 : v_dec_inst_0 = data[31:0];
	    8'b10100110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10100101 : v_dec_inst_0 = data[31:0];
	    8'b10100100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10100011 : v_dec_inst_0 = data[31:0];
	    8'b10100010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10100001 : v_dec_inst_0 = data[31:0];
	    8'b10100000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10011111 : v_dec_inst_0 = data[31:0];
	    8'b10011110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10011101 : v_dec_inst_0 = data[31:0];
	    8'b10011100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10011011 : v_dec_inst_0 = data[31:0];
	    8'b10011010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10011001 : v_dec_inst_0 = data[31:0];
	    8'b10011000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10010111 : v_dec_inst_0 = data[31:0];
	    8'b10010110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10010101 : v_dec_inst_0 = data[31:0];
	    8'b10010100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10010011 : v_dec_inst_0 = data[31:0];
	    8'b10010010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10010001 : v_dec_inst_0 = data[31:0];
	    8'b10010000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10001111 : v_dec_inst_0 = data[31:0];
	    8'b10001110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10001101 : v_dec_inst_0 = data[31:0];
	    8'b10001100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10001011 : v_dec_inst_0 = data[31:0];
	    8'b10001010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10001001 : v_dec_inst_0 = data[31:0];
	    8'b10001000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10000111 : v_dec_inst_0 = data[31:0];
	    8'b10000110 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10000101 : v_dec_inst_0 = data[31:0];
	    8'b10000100 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10000011 : v_dec_inst_0 = data[31:0];
	    8'b10000010 : v_dec_inst_0 = {16'b0, data[15:0]};
	    8'b10000001 : v_dec_inst_0 = data[31:0];
	    8'b10000000 : v_dec_inst_0 = {16'b0, data[15:0]};
	    default : v_dec_inst_0 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1111110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1111101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1111100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1111011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1111010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1111001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1111000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1110111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1110110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1110101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1110100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1110011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1110010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1110001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1110000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1101111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1101110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1101101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1101100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1101011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1101010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1101001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1101000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1100111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1100110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1100101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1100100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1100011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1100010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1100001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1100000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1011111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1011110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1011101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1011100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1011011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1011010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1011001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1011000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1010111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1010110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1010101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1010100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1010011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1010010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1010001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1010000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1001111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1001110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1001101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1001100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1001011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1001010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1001001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1001000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1000111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1000110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1000101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1000100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1000011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1000010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1000001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1000000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b111111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b111110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b111101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b111100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b111011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b111010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b111001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b111000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b110111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b110110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b110101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b110100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b110011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b110010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b110001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b110000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b101111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b101110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b101101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b101100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b101011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b101010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b101001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b101000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b100111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b100110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b100101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b100100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b100011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b100010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b100001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b100000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b1000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b1 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b0 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11111111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11111110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11111101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11111100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11111011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11111010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11111001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11111000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11110111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11110110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11110101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11110100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11110011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11110010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11110001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11110000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11101111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11101110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11101101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11101100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11101011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11101010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11101001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11101000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11100111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11100110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11100101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11100100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11100011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11100010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11100001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11100000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11011111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11011110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11011101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11011100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11011011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11011010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11011001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11011000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11010111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11010110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11010101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11010100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11010011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11010010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11010001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11010000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11001111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11001110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11001101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11001100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11001011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11001010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11001001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11001000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11000111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11000110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11000101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11000100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11000011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11000010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b11000001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b11000000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10111111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10111110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10111101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10111100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10111011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10111010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10111001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10111000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10110111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10110110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10110101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10110100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10110011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10110010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10110001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10110000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10101111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10101110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10101101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10101100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10101011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10101010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10101001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10101000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10100111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10100110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10100101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10100100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10100011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10100010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10100001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10100000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10011111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10011110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10011101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10011100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10011011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10011010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10011001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10011000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10010111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10010110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10010101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10010100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10010011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10010010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10010001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10010000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10001111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10001110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10001101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10001100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10001011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10001010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10001001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10001000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10000111 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10000110 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10000101 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10000100 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10000011 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10000010 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    8'b10000001 : v_dec_ena_0 = (v_ena[0] && v_vld[1]);
	    8'b10000000 : v_dec_ena_0 = (v_ena[0] && v_vld[0]);
	    default : v_dec_ena_0 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1111110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1111101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1111100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1111011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1111010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1111001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1111000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1110111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1110110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1110101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1110100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1110011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1110010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1110001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1110000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1101111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1101110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1101101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1101100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1101011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1101010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1101001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1101000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1100111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1100110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1100101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1100100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1100011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1100010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1100001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1100000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1011111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1011110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1011101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1011100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1011011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1011010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1011001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1011000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1010111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1010110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1010101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1010100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1010011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1010010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1010001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1010000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1001111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1001110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1001101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1001100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1001011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1001010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1001001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1001000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1000111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1000110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1000101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1000100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1000011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1000010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1000001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1000000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b111111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b111110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b111101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b111100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b111011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b111010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b111001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b111000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b110111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b110110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b110101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b110100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b110011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b110010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b110001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b110000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b101111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b101110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b101101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b101100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b101011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b101010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b101001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b101000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b100111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b100110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b100101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b100100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b100011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b100010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b100001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b100000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b1000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b1 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b0 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11111111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11111110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11111101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11111100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11111011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11111010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11111001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11111000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11110111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11110110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11110101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11110100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11110011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11110010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11110001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11110000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11101111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11101110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11101101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11101100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11101011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11101010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11101001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11101000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11100111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11100110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11100101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11100100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11100011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11100010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11100001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11100000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11011111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11011110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11011101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11011100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11011011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11011010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11011001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11011000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11010111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11010110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11010101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11010100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11010011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11010010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11010001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11010000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11001111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11001110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11001101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11001100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11001011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11001010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11001001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11001000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11000111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11000110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11000101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11000100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11000011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11000010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b11000001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b11000000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10111111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10111110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10111101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10111100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10111011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10111010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10111001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10111000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10110111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10110110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10110101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10110100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10110011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10110010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10110001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10110000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10101111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10101110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10101101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10101100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10101011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10101010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10101001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10101000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10100111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10100110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10100101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10100100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10100011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10100010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10100001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10100000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10011111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10011110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10011101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10011100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10011011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10011010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10011001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10011000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10010111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10010110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10010101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10010100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10010011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10010010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10010001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10010000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10001111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10001110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10001101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10001100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10001011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10001010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10001001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10001000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10000111 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10000110 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10000101 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10000100 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10000011 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10000010 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    8'b10000001 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[1]));
	    8'b10000000 : v_dec_vld_0 = (v_ena[0] && (v_ena[0] ^ v_vld[0]));
	    default : v_dec_vld_0 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1111110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1111101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1111100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1111011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1111010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1111001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1111000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1110111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1110110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1110101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1110100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1110011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1110010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1110001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1110000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1101111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1101110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1101101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1101100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1101011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1101010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1101001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1101000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1100111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1100110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1100101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1100100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1100011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1100010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1100001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1100000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1011111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1011110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1011101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1011100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1011011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1011010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1011001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1011000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1010111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1010110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1010101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1010100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1010011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1010010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1010001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1010000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1001111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1001110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1001101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1001100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1001011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1001010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1001001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1001000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1000111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1000110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1000101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1000100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1000011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1000010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1000001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1000000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b111111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b111110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b111101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b111100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b111011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b111010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b111001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b111000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b110111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b110110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b110101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b110100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b110011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b110010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b110001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b110000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b101111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b101110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b101101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b101100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b101011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b101010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b101001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b101000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b100111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b100110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b100101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b100100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b100011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b100010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b100001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b100000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b1000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b1 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b0 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11111111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11111110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11111101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11111100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11111011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11111010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11111001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11111000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11110111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11110110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11110101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11110100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11110011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11110010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11110001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11110000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11101111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11101110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11101101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11101100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11101011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11101010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11101001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11101000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11100111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11100110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11100101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11100100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11100011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11100010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11100001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11100000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11011111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11011110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11011101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11011100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11011011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11011010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11011001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11011000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11010111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11010110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11010101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11010100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11010011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11010010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11010001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11010000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11001111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11001110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11001101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11001100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11001011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11001010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11001001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11001000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11000111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11000110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11000101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11000100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11000011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11000010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b11000001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b11000000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10111111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10111110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10111101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10111100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10111011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10111010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10111001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10111000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10110111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10110110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10110101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10110100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10110011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10110010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10110001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10110000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10101111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10101110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10101101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10101100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10101011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10101010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10101001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10101000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10100111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10100110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10100101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10100100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10100011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10100010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10100001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10100000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10011111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10011110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10011101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10011100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10011011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10011010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10011001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10011000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10010111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10010110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10010101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10010100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10010011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10010010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10010001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10010000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10001111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10001110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10001101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10001100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10001011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10001010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10001001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10001000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10000111 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10000110 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10000101 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10000100 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10000011 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10000010 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    8'b10000001 : v_dec_pc_add_0 = (pred_pc + 32'b100);
	    8'b10000000 : v_dec_pc_add_0 = (pred_pc + 32'b10);
	    default : v_dec_pc_add_0 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_inst_1 = data[63:32];
	    8'b1111110 : v_dec_inst_1 = data[47:16];
	    8'b1111101 : v_dec_inst_1 = data[63:32];
	    8'b1111100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1111011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1111010 : v_dec_inst_1 = data[47:16];
	    8'b1111001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1111000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1110111 : v_dec_inst_1 = data[63:32];
	    8'b1110110 : v_dec_inst_1 = data[47:16];
	    8'b1110101 : v_dec_inst_1 = data[63:32];
	    8'b1110100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1110011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1110010 : v_dec_inst_1 = data[47:16];
	    8'b1110001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1110000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1101111 : v_dec_inst_1 = data[63:32];
	    8'b1101110 : v_dec_inst_1 = data[47:16];
	    8'b1101101 : v_dec_inst_1 = data[63:32];
	    8'b1101100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1101011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1101010 : v_dec_inst_1 = data[47:16];
	    8'b1101001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1101000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1100111 : v_dec_inst_1 = data[63:32];
	    8'b1100110 : v_dec_inst_1 = data[47:16];
	    8'b1100101 : v_dec_inst_1 = data[63:32];
	    8'b1100100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1100011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1100010 : v_dec_inst_1 = data[47:16];
	    8'b1100001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1100000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1011111 : v_dec_inst_1 = data[63:32];
	    8'b1011110 : v_dec_inst_1 = data[47:16];
	    8'b1011101 : v_dec_inst_1 = data[63:32];
	    8'b1011100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1011011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1011010 : v_dec_inst_1 = data[47:16];
	    8'b1011001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1011000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1010111 : v_dec_inst_1 = data[63:32];
	    8'b1010110 : v_dec_inst_1 = data[47:16];
	    8'b1010101 : v_dec_inst_1 = data[63:32];
	    8'b1010100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1010011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1010010 : v_dec_inst_1 = data[47:16];
	    8'b1010001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1010000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1001111 : v_dec_inst_1 = data[63:32];
	    8'b1001110 : v_dec_inst_1 = data[47:16];
	    8'b1001101 : v_dec_inst_1 = data[63:32];
	    8'b1001100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1001011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1001010 : v_dec_inst_1 = data[47:16];
	    8'b1001001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1001000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1000111 : v_dec_inst_1 = data[63:32];
	    8'b1000110 : v_dec_inst_1 = data[47:16];
	    8'b1000101 : v_dec_inst_1 = data[63:32];
	    8'b1000100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1000011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1000010 : v_dec_inst_1 = data[47:16];
	    8'b1000001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1000000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b111111 : v_dec_inst_1 = data[63:32];
	    8'b111110 : v_dec_inst_1 = data[47:16];
	    8'b111101 : v_dec_inst_1 = data[63:32];
	    8'b111100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b111011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b111010 : v_dec_inst_1 = data[47:16];
	    8'b111001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b111000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b110111 : v_dec_inst_1 = data[63:32];
	    8'b110110 : v_dec_inst_1 = data[47:16];
	    8'b110101 : v_dec_inst_1 = data[63:32];
	    8'b110100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b110011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b110010 : v_dec_inst_1 = data[47:16];
	    8'b110001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b110000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b101111 : v_dec_inst_1 = data[63:32];
	    8'b101110 : v_dec_inst_1 = data[47:16];
	    8'b101101 : v_dec_inst_1 = data[63:32];
	    8'b101100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b101011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b101010 : v_dec_inst_1 = data[47:16];
	    8'b101001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b101000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b100111 : v_dec_inst_1 = data[63:32];
	    8'b100110 : v_dec_inst_1 = data[47:16];
	    8'b100101 : v_dec_inst_1 = data[63:32];
	    8'b100100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b100011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b100010 : v_dec_inst_1 = data[47:16];
	    8'b100001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b100000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11111 : v_dec_inst_1 = data[63:32];
	    8'b11110 : v_dec_inst_1 = data[47:16];
	    8'b11101 : v_dec_inst_1 = data[63:32];
	    8'b11100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11010 : v_dec_inst_1 = data[47:16];
	    8'b11001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10111 : v_dec_inst_1 = data[63:32];
	    8'b10110 : v_dec_inst_1 = data[47:16];
	    8'b10101 : v_dec_inst_1 = data[63:32];
	    8'b10100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10010 : v_dec_inst_1 = data[47:16];
	    8'b10001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1111 : v_dec_inst_1 = data[63:32];
	    8'b1110 : v_dec_inst_1 = data[47:16];
	    8'b1101 : v_dec_inst_1 = data[63:32];
	    8'b1100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b1011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1010 : v_dec_inst_1 = data[47:16];
	    8'b1001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b1000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b111 : v_dec_inst_1 = data[63:32];
	    8'b110 : v_dec_inst_1 = data[47:16];
	    8'b101 : v_dec_inst_1 = data[63:32];
	    8'b100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10 : v_dec_inst_1 = data[47:16];
	    8'b1 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b0 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11111111 : v_dec_inst_1 = data[63:32];
	    8'b11111110 : v_dec_inst_1 = data[47:16];
	    8'b11111101 : v_dec_inst_1 = data[63:32];
	    8'b11111100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11111011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11111010 : v_dec_inst_1 = data[47:16];
	    8'b11111001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11111000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11110111 : v_dec_inst_1 = data[63:32];
	    8'b11110110 : v_dec_inst_1 = data[47:16];
	    8'b11110101 : v_dec_inst_1 = data[63:32];
	    8'b11110100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11110011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11110010 : v_dec_inst_1 = data[47:16];
	    8'b11110001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11110000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11101111 : v_dec_inst_1 = data[63:32];
	    8'b11101110 : v_dec_inst_1 = data[47:16];
	    8'b11101101 : v_dec_inst_1 = data[63:32];
	    8'b11101100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11101011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11101010 : v_dec_inst_1 = data[47:16];
	    8'b11101001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11101000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11100111 : v_dec_inst_1 = data[63:32];
	    8'b11100110 : v_dec_inst_1 = data[47:16];
	    8'b11100101 : v_dec_inst_1 = data[63:32];
	    8'b11100100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11100011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11100010 : v_dec_inst_1 = data[47:16];
	    8'b11100001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11100000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11011111 : v_dec_inst_1 = data[63:32];
	    8'b11011110 : v_dec_inst_1 = data[47:16];
	    8'b11011101 : v_dec_inst_1 = data[63:32];
	    8'b11011100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11011011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11011010 : v_dec_inst_1 = data[47:16];
	    8'b11011001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11011000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11010111 : v_dec_inst_1 = data[63:32];
	    8'b11010110 : v_dec_inst_1 = data[47:16];
	    8'b11010101 : v_dec_inst_1 = data[63:32];
	    8'b11010100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11010011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11010010 : v_dec_inst_1 = data[47:16];
	    8'b11010001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11010000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11001111 : v_dec_inst_1 = data[63:32];
	    8'b11001110 : v_dec_inst_1 = data[47:16];
	    8'b11001101 : v_dec_inst_1 = data[63:32];
	    8'b11001100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11001011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11001010 : v_dec_inst_1 = data[47:16];
	    8'b11001001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11001000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11000111 : v_dec_inst_1 = data[63:32];
	    8'b11000110 : v_dec_inst_1 = data[47:16];
	    8'b11000101 : v_dec_inst_1 = data[63:32];
	    8'b11000100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b11000011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11000010 : v_dec_inst_1 = data[47:16];
	    8'b11000001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b11000000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10111111 : v_dec_inst_1 = data[63:32];
	    8'b10111110 : v_dec_inst_1 = data[47:16];
	    8'b10111101 : v_dec_inst_1 = data[63:32];
	    8'b10111100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10111011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10111010 : v_dec_inst_1 = data[47:16];
	    8'b10111001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10111000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10110111 : v_dec_inst_1 = data[63:32];
	    8'b10110110 : v_dec_inst_1 = data[47:16];
	    8'b10110101 : v_dec_inst_1 = data[63:32];
	    8'b10110100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10110011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10110010 : v_dec_inst_1 = data[47:16];
	    8'b10110001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10110000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10101111 : v_dec_inst_1 = data[63:32];
	    8'b10101110 : v_dec_inst_1 = data[47:16];
	    8'b10101101 : v_dec_inst_1 = data[63:32];
	    8'b10101100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10101011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10101010 : v_dec_inst_1 = data[47:16];
	    8'b10101001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10101000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10100111 : v_dec_inst_1 = data[63:32];
	    8'b10100110 : v_dec_inst_1 = data[47:16];
	    8'b10100101 : v_dec_inst_1 = data[63:32];
	    8'b10100100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10100011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10100010 : v_dec_inst_1 = data[47:16];
	    8'b10100001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10100000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10011111 : v_dec_inst_1 = data[63:32];
	    8'b10011110 : v_dec_inst_1 = data[47:16];
	    8'b10011101 : v_dec_inst_1 = data[63:32];
	    8'b10011100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10011011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10011010 : v_dec_inst_1 = data[47:16];
	    8'b10011001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10011000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10010111 : v_dec_inst_1 = data[63:32];
	    8'b10010110 : v_dec_inst_1 = data[47:16];
	    8'b10010101 : v_dec_inst_1 = data[63:32];
	    8'b10010100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10010011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10010010 : v_dec_inst_1 = data[47:16];
	    8'b10010001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10010000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10001111 : v_dec_inst_1 = data[63:32];
	    8'b10001110 : v_dec_inst_1 = data[47:16];
	    8'b10001101 : v_dec_inst_1 = data[63:32];
	    8'b10001100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10001011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10001010 : v_dec_inst_1 = data[47:16];
	    8'b10001001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10001000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10000111 : v_dec_inst_1 = data[63:32];
	    8'b10000110 : v_dec_inst_1 = data[47:16];
	    8'b10000101 : v_dec_inst_1 = data[63:32];
	    8'b10000100 : v_dec_inst_1 = {16'b0, data[31:16]};
	    8'b10000011 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10000010 : v_dec_inst_1 = data[47:16];
	    8'b10000001 : v_dec_inst_1 = {16'b0, data[47:32]};
	    8'b10000000 : v_dec_inst_1 = {16'b0, data[31:16]};
	    default : v_dec_inst_1 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1111110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1111101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1111100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1111011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1111010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1111001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1111000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1110111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1110110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1110101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1110100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1110011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1110010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1110001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1110000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1101111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1101110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1101101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1101100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1101011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1101010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1101001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1101000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1100111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1100110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1100101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1100100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1100011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1100010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1100001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1100000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1011111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1011110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1011101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1011100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1011011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1011010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1011001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1011000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1010111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1010110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1010101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1010100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1010011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1010010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1010001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1010000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1001111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1001110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1001101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1001100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1001011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1001010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1001001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1001000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1000111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1000110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1000101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1000100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1000011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1000010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1000001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1000000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b111111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b111110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b111101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b111100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b111011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b111010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b111001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b111000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b110111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b110110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b110101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b110100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b110011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b110010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b110001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b110000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b101111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b101110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b101101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b101100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b101011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b101010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b101001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b101000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b100111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b100110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b100101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b100100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b100011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b100010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b100001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b100000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b1100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b1011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b1000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b1 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b0 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11111111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11111110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11111101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11111100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11111011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11111010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11111001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11111000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11110111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11110110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11110101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11110100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11110011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11110010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11110001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11110000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11101111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11101110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11101101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11101100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11101011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11101010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11101001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11101000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11100111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11100110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11100101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11100100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11100011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11100010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11100001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11100000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11011111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11011110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11011101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11011100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11011011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11011010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11011001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11011000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11010111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11010110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11010101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11010100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11010011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11010010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11010001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11010000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11001111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11001110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11001101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11001100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11001011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11001010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11001001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11001000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11000111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11000110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11000101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b11000100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b11000011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11000010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b11000001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b11000000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10111111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10111110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10111101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10111100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10111011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10111010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10111001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10111000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10110111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10110110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10110101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10110100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10110011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10110010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10110001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10110000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10101111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10101110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10101101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10101100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10101011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10101010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10101001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10101000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10100111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10100110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10100101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10100100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10100011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10100010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10100001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10100000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10011111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10011110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10011101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10011100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10011011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10011010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10011001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10011000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10010111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10010110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10010101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10010100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10010011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10010010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10010001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10010000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10001111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10001110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10001101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10001100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10001011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10001010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10001001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10001000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10000111 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10000110 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10000101 : v_dec_ena_1 = (v_ena[2] && v_vld[3]);
	    8'b10000100 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    8'b10000011 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10000010 : v_dec_ena_1 = (v_ena[1] && v_vld[2]);
	    8'b10000001 : v_dec_ena_1 = (v_ena[2] && v_vld[2]);
	    8'b10000000 : v_dec_ena_1 = (v_ena[1] && v_vld[1]);
	    default : v_dec_ena_1 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1111110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1111101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1111100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1111011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1111010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1111001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1111000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1110111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1110110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1110101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1110100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1110011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1110010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1110001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1110000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1101111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1101110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1101101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1101100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1101011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1101010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1101001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1101000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1100111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1100110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1100101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1100100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1100011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1100010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1100001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1100000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1011111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1011110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1011101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1011100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1011011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1011010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1011001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1011000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1010111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1010110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1010101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1010100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1010011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1010010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1010001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1010000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1001111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1001110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1001101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1001100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1001011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1001010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1001001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1001000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1000111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1000110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1000101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1000100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1000011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1000010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1000001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1000000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b111111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b111110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b111101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b111100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b111011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b111010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b111001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b111000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b110111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b110110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b110101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b110100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b110011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b110010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b110001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b110000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b101111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b101110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b101101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b101100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b101011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b101010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b101001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b101000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b100111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b100110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b100101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b100100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b100011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b100010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b100001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b100000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b1011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b1 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b0 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11111111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11111110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11111101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11111100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11111011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11111010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11111001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11111000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11110111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11110110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11110101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11110100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11110011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11110010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11110001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11110000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11101111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11101110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11101101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11101100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11101011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11101010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11101001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11101000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11100111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11100110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11100101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11100100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11100011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11100010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11100001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11100000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11011111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11011110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11011101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11011100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11011011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11011010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11011001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11011000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11010111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11010110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11010101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11010100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11010011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11010010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11010001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11010000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11001111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11001110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11001101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11001100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11001011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11001010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11001001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11001000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11000111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11000110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11000101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11000100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b11000011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11000010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b11000001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11000000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10111111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10111110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10111101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10111100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10111011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10111010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10111001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10111000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10110111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10110110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10110101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10110100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10110011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10110010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10110001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10110000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10101111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10101110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10101101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10101100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10101011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10101010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10101001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10101000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10100111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10100110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10100101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10100100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10100011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10100010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10100001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10100000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10011111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10011110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10011101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10011100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10011011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10011010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10011001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10011000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10010111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10010110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10010101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10010100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10010011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10010010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10010001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10010000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10001111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10001110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10001101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10001100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10001011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10001010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10001001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10001000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10000111 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10000110 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10000101 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10000100 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    8'b10000011 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10000010 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[2]));
	    8'b10000001 : v_dec_vld_1 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10000000 : v_dec_vld_1 = (v_ena[1] && (v_ena[1] ^ v_vld[1]));
	    default : v_dec_vld_1 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1111110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1111101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1111100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1111011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1111010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1111001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1111000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1110111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1110110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1110101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1110100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1110011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1110010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1110001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1110000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1101111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1101110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1101101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1101100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1101011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1101010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1101001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1101000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1100111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1100110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1100101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1100100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1100011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1100010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1100001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1100000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1011111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1011110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1011101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1011100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1011011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1011010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1011001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1011000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1010111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1010110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1010101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1010100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1010011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1010010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1010001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1010000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1001111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1001110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1001101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1001100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1001011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1001010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1001001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1001000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1000111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1000110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1000101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1000100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1000011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1000010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1000001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1000000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b111111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b111110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b111101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b111100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b111011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b111010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b111001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b111000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b110111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b110110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b110101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b110100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b110011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b110010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b110001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b110000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b101111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b101110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b101101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b101100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b101011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b101010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b101001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b101000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b100111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b100110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b100101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b100100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b100011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b100010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b100001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b100000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b1100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b1011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b1 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b0 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11111111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11111110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11111101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11111100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11111011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11111010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11111001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11111000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11110111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11110110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11110101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11110100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11110011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11110010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11110001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11110000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11101111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11101110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11101101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11101100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11101011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11101010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11101001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11101000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11100111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11100110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11100101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11100100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11100011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11100010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11100001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11100000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11011111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11011110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11011101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11011100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11011011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11011010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11011001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11011000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11010111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11010110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11010101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11010100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11010011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11010010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11010001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11010000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11001111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11001110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11001101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11001100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11001011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11001010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11001001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11001000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11000111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11000110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11000101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b11000100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b11000011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11000010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11000001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b11000000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10111111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10111110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10111101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10111100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10111011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10111010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10111001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10111000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10110111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10110110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10110101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10110100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10110011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10110010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10110001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10110000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10101111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10101110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10101101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10101100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10101011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10101010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10101001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10101000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10100111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10100110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10100101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10100100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10100011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10100010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10100001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10100000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10011111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10011110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10011101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10011100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10011011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10011010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10011001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10011000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10010111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10010110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10010101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10010100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10010011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10010010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10010001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10010000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10001111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10001110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10001101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10001100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10001011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10001010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10001001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10001000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10000111 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10000110 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10000101 : v_dec_pc_add_1 = (pred_pc + 32'b1000);
	    8'b10000100 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    8'b10000011 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10000010 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10000001 : v_dec_pc_add_1 = (pred_pc + 32'b110);
	    8'b10000000 : v_dec_pc_add_1 = (pred_pc + 32'b100);
	    default : v_dec_pc_add_1 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_inst_2 = data[95:64];
	    8'b1111110 : v_dec_inst_2 = data[79:48];
	    8'b1111101 : v_dec_inst_2 = data[95:64];
	    8'b1111100 : v_dec_inst_2 = data[63:32];
	    8'b1111011 : v_dec_inst_2 = data[79:48];
	    8'b1111010 : v_dec_inst_2 = data[79:48];
	    8'b1111001 : v_dec_inst_2 = data[79:48];
	    8'b1111000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1110111 : v_dec_inst_2 = data[95:64];
	    8'b1110110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1110101 : v_dec_inst_2 = data[95:64];
	    8'b1110100 : v_dec_inst_2 = data[63:32];
	    8'b1110011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1110010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1110001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1110000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1101111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1101110 : v_dec_inst_2 = data[79:48];
	    8'b1101101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1101100 : v_dec_inst_2 = data[63:32];
	    8'b1101011 : v_dec_inst_2 = data[79:48];
	    8'b1101010 : v_dec_inst_2 = data[79:48];
	    8'b1101001 : v_dec_inst_2 = data[79:48];
	    8'b1101000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1100111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1100110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1100101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1100100 : v_dec_inst_2 = data[63:32];
	    8'b1100011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1100010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1100001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1100000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1011111 : v_dec_inst_2 = data[95:64];
	    8'b1011110 : v_dec_inst_2 = data[79:48];
	    8'b1011101 : v_dec_inst_2 = data[95:64];
	    8'b1011100 : v_dec_inst_2 = data[63:32];
	    8'b1011011 : v_dec_inst_2 = data[79:48];
	    8'b1011010 : v_dec_inst_2 = data[79:48];
	    8'b1011001 : v_dec_inst_2 = data[79:48];
	    8'b1011000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1010111 : v_dec_inst_2 = data[95:64];
	    8'b1010110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1010101 : v_dec_inst_2 = data[95:64];
	    8'b1010100 : v_dec_inst_2 = data[63:32];
	    8'b1010011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1010010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1010001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1010000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1001111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1001110 : v_dec_inst_2 = data[79:48];
	    8'b1001101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1001100 : v_dec_inst_2 = data[63:32];
	    8'b1001011 : v_dec_inst_2 = data[79:48];
	    8'b1001010 : v_dec_inst_2 = data[79:48];
	    8'b1001001 : v_dec_inst_2 = data[79:48];
	    8'b1001000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1000111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1000110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1000101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1000100 : v_dec_inst_2 = data[63:32];
	    8'b1000011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1000010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1000001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1000000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b111111 : v_dec_inst_2 = data[95:64];
	    8'b111110 : v_dec_inst_2 = data[79:48];
	    8'b111101 : v_dec_inst_2 = data[95:64];
	    8'b111100 : v_dec_inst_2 = data[63:32];
	    8'b111011 : v_dec_inst_2 = data[79:48];
	    8'b111010 : v_dec_inst_2 = data[79:48];
	    8'b111001 : v_dec_inst_2 = data[79:48];
	    8'b111000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b110111 : v_dec_inst_2 = data[95:64];
	    8'b110110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b110101 : v_dec_inst_2 = data[95:64];
	    8'b110100 : v_dec_inst_2 = data[63:32];
	    8'b110011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b110010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b110001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b110000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b101111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b101110 : v_dec_inst_2 = data[79:48];
	    8'b101101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b101100 : v_dec_inst_2 = data[63:32];
	    8'b101011 : v_dec_inst_2 = data[79:48];
	    8'b101010 : v_dec_inst_2 = data[79:48];
	    8'b101001 : v_dec_inst_2 = data[79:48];
	    8'b101000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b100111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b100110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b100101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b100100 : v_dec_inst_2 = data[63:32];
	    8'b100011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b100010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b100001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b100000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11111 : v_dec_inst_2 = data[95:64];
	    8'b11110 : v_dec_inst_2 = data[79:48];
	    8'b11101 : v_dec_inst_2 = data[95:64];
	    8'b11100 : v_dec_inst_2 = data[63:32];
	    8'b11011 : v_dec_inst_2 = data[79:48];
	    8'b11010 : v_dec_inst_2 = data[79:48];
	    8'b11001 : v_dec_inst_2 = data[79:48];
	    8'b11000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10111 : v_dec_inst_2 = data[95:64];
	    8'b10110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10101 : v_dec_inst_2 = data[95:64];
	    8'b10100 : v_dec_inst_2 = data[63:32];
	    8'b10011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b1111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1110 : v_dec_inst_2 = data[79:48];
	    8'b1101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b1100 : v_dec_inst_2 = data[63:32];
	    8'b1011 : v_dec_inst_2 = data[79:48];
	    8'b1010 : v_dec_inst_2 = data[79:48];
	    8'b1001 : v_dec_inst_2 = data[79:48];
	    8'b1000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b100 : v_dec_inst_2 = data[63:32];
	    8'b11 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b1 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b0 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11111111 : v_dec_inst_2 = data[95:64];
	    8'b11111110 : v_dec_inst_2 = data[79:48];
	    8'b11111101 : v_dec_inst_2 = data[95:64];
	    8'b11111100 : v_dec_inst_2 = data[63:32];
	    8'b11111011 : v_dec_inst_2 = data[79:48];
	    8'b11111010 : v_dec_inst_2 = data[79:48];
	    8'b11111001 : v_dec_inst_2 = data[79:48];
	    8'b11111000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11110111 : v_dec_inst_2 = data[95:64];
	    8'b11110110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11110101 : v_dec_inst_2 = data[95:64];
	    8'b11110100 : v_dec_inst_2 = data[63:32];
	    8'b11110011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11110010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11110001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11110000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11101111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11101110 : v_dec_inst_2 = data[79:48];
	    8'b11101101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11101100 : v_dec_inst_2 = data[63:32];
	    8'b11101011 : v_dec_inst_2 = data[79:48];
	    8'b11101010 : v_dec_inst_2 = data[79:48];
	    8'b11101001 : v_dec_inst_2 = data[79:48];
	    8'b11101000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11100111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11100110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11100101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11100100 : v_dec_inst_2 = data[63:32];
	    8'b11100011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11100010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11100001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11100000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11011111 : v_dec_inst_2 = data[95:64];
	    8'b11011110 : v_dec_inst_2 = data[79:48];
	    8'b11011101 : v_dec_inst_2 = data[95:64];
	    8'b11011100 : v_dec_inst_2 = data[63:32];
	    8'b11011011 : v_dec_inst_2 = data[79:48];
	    8'b11011010 : v_dec_inst_2 = data[79:48];
	    8'b11011001 : v_dec_inst_2 = data[79:48];
	    8'b11011000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11010111 : v_dec_inst_2 = data[95:64];
	    8'b11010110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11010101 : v_dec_inst_2 = data[95:64];
	    8'b11010100 : v_dec_inst_2 = data[63:32];
	    8'b11010011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11010010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11010001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11010000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11001111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11001110 : v_dec_inst_2 = data[79:48];
	    8'b11001101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11001100 : v_dec_inst_2 = data[63:32];
	    8'b11001011 : v_dec_inst_2 = data[79:48];
	    8'b11001010 : v_dec_inst_2 = data[79:48];
	    8'b11001001 : v_dec_inst_2 = data[79:48];
	    8'b11001000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b11000111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11000110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11000101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b11000100 : v_dec_inst_2 = data[63:32];
	    8'b11000011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11000010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11000001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b11000000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10111111 : v_dec_inst_2 = data[95:64];
	    8'b10111110 : v_dec_inst_2 = data[79:48];
	    8'b10111101 : v_dec_inst_2 = data[95:64];
	    8'b10111100 : v_dec_inst_2 = data[63:32];
	    8'b10111011 : v_dec_inst_2 = data[79:48];
	    8'b10111010 : v_dec_inst_2 = data[79:48];
	    8'b10111001 : v_dec_inst_2 = data[79:48];
	    8'b10111000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10110111 : v_dec_inst_2 = data[95:64];
	    8'b10110110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10110101 : v_dec_inst_2 = data[95:64];
	    8'b10110100 : v_dec_inst_2 = data[63:32];
	    8'b10110011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10110010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10110001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10110000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10101111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10101110 : v_dec_inst_2 = data[79:48];
	    8'b10101101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10101100 : v_dec_inst_2 = data[63:32];
	    8'b10101011 : v_dec_inst_2 = data[79:48];
	    8'b10101010 : v_dec_inst_2 = data[79:48];
	    8'b10101001 : v_dec_inst_2 = data[79:48];
	    8'b10101000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10100111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10100110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10100101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10100100 : v_dec_inst_2 = data[63:32];
	    8'b10100011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10100010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10100001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10100000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10011111 : v_dec_inst_2 = data[95:64];
	    8'b10011110 : v_dec_inst_2 = data[79:48];
	    8'b10011101 : v_dec_inst_2 = data[95:64];
	    8'b10011100 : v_dec_inst_2 = data[63:32];
	    8'b10011011 : v_dec_inst_2 = data[79:48];
	    8'b10011010 : v_dec_inst_2 = data[79:48];
	    8'b10011001 : v_dec_inst_2 = data[79:48];
	    8'b10011000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10010111 : v_dec_inst_2 = data[95:64];
	    8'b10010110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10010101 : v_dec_inst_2 = data[95:64];
	    8'b10010100 : v_dec_inst_2 = data[63:32];
	    8'b10010011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10010010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10010001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10010000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10001111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10001110 : v_dec_inst_2 = data[79:48];
	    8'b10001101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10001100 : v_dec_inst_2 = data[63:32];
	    8'b10001011 : v_dec_inst_2 = data[79:48];
	    8'b10001010 : v_dec_inst_2 = data[79:48];
	    8'b10001001 : v_dec_inst_2 = data[79:48];
	    8'b10001000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    8'b10000111 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10000110 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10000101 : v_dec_inst_2 = {16'b0, data[79:64]};
	    8'b10000100 : v_dec_inst_2 = data[63:32];
	    8'b10000011 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10000010 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10000001 : v_dec_inst_2 = {16'b0, data[63:48]};
	    8'b10000000 : v_dec_inst_2 = {16'b0, data[47:32]};
	    default : v_dec_inst_2 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1111110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1111101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1111100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1111011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1111010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1111001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1111000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1110111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1110110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1110101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1110100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1110011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1110010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1110001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1110000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1101111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1101110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1101101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1101100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1101011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1101010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1101001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1101000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1100111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1100110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1100101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1100100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1100011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1100010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1100001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1100000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1011111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1011110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1011101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1011100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1011011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1011010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1011001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1011000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1010111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1010110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1010101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b1010100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1010011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1010010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1010001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1010000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1001111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1001110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1001101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1001100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1001011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1001010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1001001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1001000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1000111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1000110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1000101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1000100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1000011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1000010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1000001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1000000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b111111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b111110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b111101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b111100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b111011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b111010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b111001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b111000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b110111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b110110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b110101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b110100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b110011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b110010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b110001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b110000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b101111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b101110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b101101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b101100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b101011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b101010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b101001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b101000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b100111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b100110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b100101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b100100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b100011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b100010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b100001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b100000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b1111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b1100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b1011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b1000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b1 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b0 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11111111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11111110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11111101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11111100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11111011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11111010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11111001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11111000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11110111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11110110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11110101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11110100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11110011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11110010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11110001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11110000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11101111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11101110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11101101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11101100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11101011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11101010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11101001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11101000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11100111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11100110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11100101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11100100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11100011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11100010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11100001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11100000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11011111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11011110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11011101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11011100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11011011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11011010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11011001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11011000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11010111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11010110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11010101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b11010100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11010011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11010010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11010001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11010000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11001111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11001110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11001101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11001100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11001011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11001010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11001001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b11001000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b11000111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11000110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11000101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b11000100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b11000011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11000010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11000001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b11000000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10111111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10111110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10111101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10111100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10111011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10111010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10111001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10111000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10110111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10110110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10110101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10110100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10110011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10110010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10110001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10110000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10101111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10101110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10101101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10101100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10101011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10101010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10101001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10101000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10100111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10100110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10100101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10100100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10100011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10100010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10100001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10100000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10011111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10011110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10011101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10011100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10011011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10011010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10011001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10011000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10010111 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10010110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10010101 : v_dec_ena_2 = (v_ena[4] && v_vld[5]);
	    8'b10010100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10010011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10010010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10010001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10010000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10001111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10001110 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10001101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10001100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10001011 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10001010 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10001001 : v_dec_ena_2 = (v_ena[3] && v_vld[4]);
	    8'b10001000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    8'b10000111 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10000110 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10000101 : v_dec_ena_2 = (v_ena[4] && v_vld[4]);
	    8'b10000100 : v_dec_ena_2 = (v_ena[2] && v_vld[3]);
	    8'b10000011 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10000010 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10000001 : v_dec_ena_2 = (v_ena[3] && v_vld[3]);
	    8'b10000000 : v_dec_ena_2 = (v_ena[2] && v_vld[2]);
	    default : v_dec_ena_2 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1111110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1111101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1111100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1111011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1111010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1111001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1111000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1110111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1110101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1110011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1110010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1110001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1110000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1101111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1101110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1101101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1101100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1101011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1101010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1101001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1101000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1100111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1100101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1100011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1100010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1100001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1100000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1011111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1011110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1011101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1011100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1011011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1011010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1011001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1011000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1010111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1010101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1010011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1010010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1010001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1010000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1001111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1001110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1001101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1001100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1001011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1001010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1001001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1001000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1000111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1000101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1000011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1000010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1000001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1000000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b111111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b111110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b111101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b111100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b111011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b111010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b111001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b111000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b110111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b110101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b110011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b110010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b110001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b110000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b101111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b101110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b101101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b101100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b101011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b101010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b101001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b101000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b100111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b100101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b100011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b100010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b100001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b100000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b1111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b1011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b0 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11111111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11111110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11111101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11111100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11111011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11111010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11111001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11111000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11110111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11110101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11110011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11110010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11110001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11110000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11101111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11101110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11101101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11101100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11101011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11101010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11101001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11101000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11100111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11100101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11100011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11100010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11100001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11100000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11011111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11011110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11011101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11011100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11011011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11011010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11011001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11011000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11010111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11010101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11010011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11010010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11010001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11010000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11001111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11001110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11001101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11001100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11001011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11001010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11001001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11001000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b11000111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11000101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b11000011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11000010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11000001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11000000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10111111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10111110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10111101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10111100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10111011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10111010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10111001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10111000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10110111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10110101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10110011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10110010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10110001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10110000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10101111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10101110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10101101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10101100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10101011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10101010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10101001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10101000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10100111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10100101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10100011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10100010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10100001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10100000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10011111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10011110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10011101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10011100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10011011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10011010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10011001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10011000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10010111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10010101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10010011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10010010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10010001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10010000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10001111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10001110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10001101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10001100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10001011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10001010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10001001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10001000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    8'b10000111 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000110 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10000101 : v_dec_vld_2 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000100 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[3]));
	    8'b10000011 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10000010 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10000001 : v_dec_vld_2 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10000000 : v_dec_vld_2 = (v_ena[2] && (v_ena[2] ^ v_vld[2]));
	    default : v_dec_vld_2 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1111110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1111101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1111100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1111011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1111010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1111001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1111000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1110111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1110110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1110101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1110100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1110011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1110010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1110001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1110000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1101111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1101011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1100111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1100110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1100101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1100100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1100011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1100010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1100001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1100000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1011111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1011110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1011101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1011100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1011011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1011010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1011001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1011000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1010111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1010110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1010101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b1010100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1010011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1010010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1010001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1010000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1001111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1001011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1000111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1000110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1000101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1000100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1000011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1000010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1000001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1000000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b111111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b111110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b111101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b111100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b111011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b111010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b111001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b111000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b110111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b110110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b110101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b110100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b110011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b110010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b110001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b110000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b101111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b101011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b101000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b100111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b100110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b100101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b100100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b100011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b100010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b100001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b100000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b1111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b1000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b1 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b0 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11111111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11111110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11111101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11111100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11111011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11111010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11111001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11111000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11110111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11110110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11110101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11110100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11110011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11110010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11110001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11110000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11101111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11101011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11101000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11100111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11100110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11100101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11100100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11100011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11100010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11100001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11100000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11011111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11011110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11011101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11011100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11011011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11011010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11011001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11011000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11010111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11010110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11010101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b11010100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11010011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11010010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11010001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11010000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11001111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11001011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11001000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b11000111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11000110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11000101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b11000100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11000011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11000010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11000001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b11000000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10111111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10111110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10111101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10111100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10111011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10111010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10111001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10111000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10110111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10110110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10110101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10110100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10110011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10110010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10110001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10110000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10101111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10101011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10101000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10100111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10100110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10100101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10100100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10100011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10100010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10100001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10100000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10011111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10011110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10011101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10011100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10011011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10011010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10011001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10011000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10010111 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10010110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010101 : v_dec_pc_add_2 = (pred_pc + 32'b1100);
	    8'b10010100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10010000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10001111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001110 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10001011 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001010 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001001 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10001000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    8'b10000111 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10000110 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000101 : v_dec_pc_add_2 = (pred_pc + 32'b1010);
	    8'b10000100 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000011 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000010 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000001 : v_dec_pc_add_2 = (pred_pc + 32'b1000);
	    8'b10000000 : v_dec_pc_add_2 = (pred_pc + 32'b110);
	    default : v_dec_pc_add_2 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_inst_3 = data[127:96];
	    8'b1111110 : v_dec_inst_3 = data[111:80];
	    8'b1111101 : v_dec_inst_3 = data[127:96];
	    8'b1111100 : v_dec_inst_3 = data[95:64];
	    8'b1111011 : v_dec_inst_3 = data[111:80];
	    8'b1111010 : v_dec_inst_3 = data[111:80];
	    8'b1111001 : v_dec_inst_3 = data[111:80];
	    8'b1111000 : v_dec_inst_3 = data[79:48];
	    8'b1110111 : v_dec_inst_3 = data[127:96];
	    8'b1110110 : v_dec_inst_3 = data[95:64];
	    8'b1110101 : v_dec_inst_3 = data[127:96];
	    8'b1110100 : v_dec_inst_3 = data[95:64];
	    8'b1110011 : v_dec_inst_3 = data[95:64];
	    8'b1110010 : v_dec_inst_3 = data[95:64];
	    8'b1110001 : v_dec_inst_3 = data[95:64];
	    8'b1110000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b1101111 : v_dec_inst_3 = data[111:80];
	    8'b1101110 : v_dec_inst_3 = data[111:80];
	    8'b1101101 : v_dec_inst_3 = data[111:80];
	    8'b1101100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1101011 : v_dec_inst_3 = data[111:80];
	    8'b1101010 : v_dec_inst_3 = data[111:80];
	    8'b1101001 : v_dec_inst_3 = data[111:80];
	    8'b1101000 : v_dec_inst_3 = data[79:48];
	    8'b1100111 : v_dec_inst_3 = data[111:80];
	    8'b1100110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1100101 : v_dec_inst_3 = data[111:80];
	    8'b1100100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1100011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1100010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1100001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1100000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b1011111 : v_dec_inst_3 = data[127:96];
	    8'b1011110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1011101 : v_dec_inst_3 = data[127:96];
	    8'b1011100 : v_dec_inst_3 = data[95:64];
	    8'b1011011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1011010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1011001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1011000 : v_dec_inst_3 = data[79:48];
	    8'b1010111 : v_dec_inst_3 = data[127:96];
	    8'b1010110 : v_dec_inst_3 = data[95:64];
	    8'b1010101 : v_dec_inst_3 = data[127:96];
	    8'b1010100 : v_dec_inst_3 = data[95:64];
	    8'b1010011 : v_dec_inst_3 = data[95:64];
	    8'b1010010 : v_dec_inst_3 = data[95:64];
	    8'b1010001 : v_dec_inst_3 = data[95:64];
	    8'b1010000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b1001111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1001011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001000 : v_dec_inst_3 = data[79:48];
	    8'b1000111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1000110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1000101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1000100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1000011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1000010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1000001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1000000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b111111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b111110 : v_dec_inst_3 = data[111:80];
	    8'b111101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b111100 : v_dec_inst_3 = data[95:64];
	    8'b111011 : v_dec_inst_3 = data[111:80];
	    8'b111010 : v_dec_inst_3 = data[111:80];
	    8'b111001 : v_dec_inst_3 = data[111:80];
	    8'b111000 : v_dec_inst_3 = data[79:48];
	    8'b110111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b110110 : v_dec_inst_3 = data[95:64];
	    8'b110101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b110100 : v_dec_inst_3 = data[95:64];
	    8'b110011 : v_dec_inst_3 = data[95:64];
	    8'b110010 : v_dec_inst_3 = data[95:64];
	    8'b110001 : v_dec_inst_3 = data[95:64];
	    8'b110000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b101111 : v_dec_inst_3 = data[111:80];
	    8'b101110 : v_dec_inst_3 = data[111:80];
	    8'b101101 : v_dec_inst_3 = data[111:80];
	    8'b101100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b101011 : v_dec_inst_3 = data[111:80];
	    8'b101010 : v_dec_inst_3 = data[111:80];
	    8'b101001 : v_dec_inst_3 = data[111:80];
	    8'b101000 : v_dec_inst_3 = data[79:48];
	    8'b100111 : v_dec_inst_3 = data[111:80];
	    8'b100110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b100101 : v_dec_inst_3 = data[111:80];
	    8'b100100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b100011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b100010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b100001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b100000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b11111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b11110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b11100 : v_dec_inst_3 = data[95:64];
	    8'b11011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11000 : v_dec_inst_3 = data[79:48];
	    8'b10111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10110 : v_dec_inst_3 = data[95:64];
	    8'b10101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10100 : v_dec_inst_3 = data[95:64];
	    8'b10011 : v_dec_inst_3 = data[95:64];
	    8'b10010 : v_dec_inst_3 = data[95:64];
	    8'b10001 : v_dec_inst_3 = data[95:64];
	    8'b10000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b1111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b1000 : v_dec_inst_3 = data[79:48];
	    8'b111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b1 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b0 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b11111111 : v_dec_inst_3 = data[127:96];
	    8'b11111110 : v_dec_inst_3 = data[111:80];
	    8'b11111101 : v_dec_inst_3 = data[127:96];
	    8'b11111100 : v_dec_inst_3 = data[95:64];
	    8'b11111011 : v_dec_inst_3 = data[111:80];
	    8'b11111010 : v_dec_inst_3 = data[111:80];
	    8'b11111001 : v_dec_inst_3 = data[111:80];
	    8'b11111000 : v_dec_inst_3 = data[79:48];
	    8'b11110111 : v_dec_inst_3 = data[127:96];
	    8'b11110110 : v_dec_inst_3 = data[95:64];
	    8'b11110101 : v_dec_inst_3 = data[127:96];
	    8'b11110100 : v_dec_inst_3 = data[95:64];
	    8'b11110011 : v_dec_inst_3 = data[95:64];
	    8'b11110010 : v_dec_inst_3 = data[95:64];
	    8'b11110001 : v_dec_inst_3 = data[95:64];
	    8'b11110000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b11101111 : v_dec_inst_3 = data[111:80];
	    8'b11101110 : v_dec_inst_3 = data[111:80];
	    8'b11101101 : v_dec_inst_3 = data[111:80];
	    8'b11101100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11101011 : v_dec_inst_3 = data[111:80];
	    8'b11101010 : v_dec_inst_3 = data[111:80];
	    8'b11101001 : v_dec_inst_3 = data[111:80];
	    8'b11101000 : v_dec_inst_3 = data[79:48];
	    8'b11100111 : v_dec_inst_3 = data[111:80];
	    8'b11100110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11100101 : v_dec_inst_3 = data[111:80];
	    8'b11100100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11100011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11100010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11100001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11100000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b11011111 : v_dec_inst_3 = data[127:96];
	    8'b11011110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11011101 : v_dec_inst_3 = data[127:96];
	    8'b11011100 : v_dec_inst_3 = data[95:64];
	    8'b11011011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11011010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11011001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11011000 : v_dec_inst_3 = data[79:48];
	    8'b11010111 : v_dec_inst_3 = data[127:96];
	    8'b11010110 : v_dec_inst_3 = data[95:64];
	    8'b11010101 : v_dec_inst_3 = data[127:96];
	    8'b11010100 : v_dec_inst_3 = data[95:64];
	    8'b11010011 : v_dec_inst_3 = data[95:64];
	    8'b11010010 : v_dec_inst_3 = data[95:64];
	    8'b11010001 : v_dec_inst_3 = data[95:64];
	    8'b11010000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b11001111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11001011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11001000 : v_dec_inst_3 = data[79:48];
	    8'b11000111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11000110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11000101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b11000100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11000011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11000010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11000001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b11000000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b10111111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10111110 : v_dec_inst_3 = data[111:80];
	    8'b10111101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10111100 : v_dec_inst_3 = data[95:64];
	    8'b10111011 : v_dec_inst_3 = data[111:80];
	    8'b10111010 : v_dec_inst_3 = data[111:80];
	    8'b10111001 : v_dec_inst_3 = data[111:80];
	    8'b10111000 : v_dec_inst_3 = data[79:48];
	    8'b10110111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10110110 : v_dec_inst_3 = data[95:64];
	    8'b10110101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10110100 : v_dec_inst_3 = data[95:64];
	    8'b10110011 : v_dec_inst_3 = data[95:64];
	    8'b10110010 : v_dec_inst_3 = data[95:64];
	    8'b10110001 : v_dec_inst_3 = data[95:64];
	    8'b10110000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b10101111 : v_dec_inst_3 = data[111:80];
	    8'b10101110 : v_dec_inst_3 = data[111:80];
	    8'b10101101 : v_dec_inst_3 = data[111:80];
	    8'b10101100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10101011 : v_dec_inst_3 = data[111:80];
	    8'b10101010 : v_dec_inst_3 = data[111:80];
	    8'b10101001 : v_dec_inst_3 = data[111:80];
	    8'b10101000 : v_dec_inst_3 = data[79:48];
	    8'b10100111 : v_dec_inst_3 = data[111:80];
	    8'b10100110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10100101 : v_dec_inst_3 = data[111:80];
	    8'b10100100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10100011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10100010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10100001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10100000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b10011111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10011110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10011101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10011100 : v_dec_inst_3 = data[95:64];
	    8'b10011011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10011010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10011001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10011000 : v_dec_inst_3 = data[79:48];
	    8'b10010111 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10010110 : v_dec_inst_3 = data[95:64];
	    8'b10010101 : v_dec_inst_3 = {16'b0, data[111:96]};
	    8'b10010100 : v_dec_inst_3 = data[95:64];
	    8'b10010011 : v_dec_inst_3 = data[95:64];
	    8'b10010010 : v_dec_inst_3 = data[95:64];
	    8'b10010001 : v_dec_inst_3 = data[95:64];
	    8'b10010000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    8'b10001111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001110 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10001011 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001010 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001001 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10001000 : v_dec_inst_3 = data[79:48];
	    8'b10000111 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10000110 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10000101 : v_dec_inst_3 = {16'b0, data[95:80]};
	    8'b10000100 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10000011 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10000010 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10000001 : v_dec_inst_3 = {16'b0, data[79:64]};
	    8'b10000000 : v_dec_inst_3 = {16'b0, data[63:48]};
	    default : v_dec_inst_3 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1111110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1111101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1111100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1111011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1111010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1111001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1111000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b1110111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1110110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1110101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1110100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1110011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1110010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1110001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1110000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b1101111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1101011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1101000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b1100111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1100110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1100101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b1100100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1100011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1100010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1100001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1100000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b1011111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1011110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1011101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1011100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1011011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1011010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1011001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1011000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b1010111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1010110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1010101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b1010100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1010011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1010010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1010001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b1010000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b1001111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1001011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b1000111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1000110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1000101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1000100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1000011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1000010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1000001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1000000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b111111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b111110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b111101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b111100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b111011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b111010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b111001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b111000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b110111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b110110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b110101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b110100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b110011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b110010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b110001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b110000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b101111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b101011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b101000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b100111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b100110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b100101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b100100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b100011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b100010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b100001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b100000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b11111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b11110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b11100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b10111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b1111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b1000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b1 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b0 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b11111111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11111110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11111101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11111100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11111011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11111010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11111001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11111000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b11110111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11110110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11110101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11110100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11110011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11110010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11110001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11110000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b11101111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11101011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11101000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b11100111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11100110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11100101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b11100100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11100011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11100010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11100001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11100000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b11011111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11011110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11011101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11011100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11011011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11011010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11011001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11011000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b11010111 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11010110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11010101 : v_dec_ena_3 = (v_ena[6] && v_vld[7]);
	    8'b11010100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11010011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11010010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11010001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b11010000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b11001111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11001011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11001000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b11000111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11000110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11000101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b11000100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11000011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11000010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11000001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b11000000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b10111111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10111110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10111101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10111100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10111011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10111010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10111001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10111000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b10110111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10110110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10110101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10110100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10110011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10110010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10110001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10110000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b10101111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101110 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10101011 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101010 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101001 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10101000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b10100111 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10100110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10100101 : v_dec_ena_3 = (v_ena[5] && v_vld[6]);
	    8'b10100100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10100011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10100010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10100001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10100000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b10011111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10011110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10011101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10011100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10011011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10011010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10011001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10011000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b10010111 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10010110 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010101 : v_dec_ena_3 = (v_ena[6] && v_vld[6]);
	    8'b10010100 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010011 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010010 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010001 : v_dec_ena_3 = (v_ena[4] && v_vld[5]);
	    8'b10010000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    8'b10001111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001110 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10001011 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001010 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001001 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10001000 : v_dec_ena_3 = (v_ena[3] && v_vld[4]);
	    8'b10000111 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10000110 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10000101 : v_dec_ena_3 = (v_ena[5] && v_vld[5]);
	    8'b10000100 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10000011 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10000010 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10000001 : v_dec_ena_3 = (v_ena[4] && v_vld[4]);
	    8'b10000000 : v_dec_ena_3 = (v_ena[3] && v_vld[3]);
	    default : v_dec_ena_3 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1111110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1111101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1111100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1111011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1111010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1111001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1111000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1110111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1110000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1101111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1101011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1100111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1100000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1011111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1011101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1011011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1011010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1011001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1011000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1010111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1010000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1001111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1001011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b1000111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1000000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b111111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b111110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b111101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b111100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b111011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b111010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b111001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b111000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b110111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b110000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b101111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b101011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b100111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b100000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b1111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b0 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11111111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11111110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11111101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11111100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11111011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11111010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11111001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11111000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11110111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11110000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11101111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11101011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11100111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11100000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11011111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11011101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11011011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11011010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11011001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11011000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11010111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11010000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b11001111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11001011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b11000111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11000000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10111111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10111110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10111101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10111100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10111011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10111010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10111001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10111000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10110111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10110000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10101111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10101011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10100111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10100000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10011111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10011101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10011011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10011010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10011001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10011000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10010111 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010101 : v_dec_vld_3 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10010000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    8'b10001111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001110 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10001011 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001010 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001001 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[4]));
	    8'b10000111 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000110 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000101 : v_dec_vld_3 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000100 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000011 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000010 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000001 : v_dec_vld_3 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10000000 : v_dec_vld_3 = (v_ena[3] && (v_ena[3] ^ v_vld[3]));
	    default : v_dec_vld_3 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1111110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1111101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1111100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1111011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1111010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1111001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1111000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1110111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1110110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1110100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b1101111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1101011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1101000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1100110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b1100100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1100000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b1011111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1011110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1011101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1011100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1011011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1011010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1011001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1011000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1010111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1010110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b1010100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b1001111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1001011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1000110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1000100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1000000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b111111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b111011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b111000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b110111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b110110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b110100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b101111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b101011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b101000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b100110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b100100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b100000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b11111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b1111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b1000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b1 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b0 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b11111111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11111110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11111101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11111100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11111011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11111010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11111001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11111000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11110111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11110110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11110101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11110100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11110011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11110010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11110001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11110000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b11101111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11101011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11101000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11100110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b11100100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11100000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b11011111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11011110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11011100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11011000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11010111 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11010110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010101 : v_dec_pc_add_3 = (pred_pc + 32'b10000);
	    8'b11010100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11010000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b11001111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11001011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11001000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11000110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b11000100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b11000000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b10111111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10111011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10111000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10110111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10110110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10110101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10110100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10110011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10110010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10110001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10110000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b10101111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101110 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10101011 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101010 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101001 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10101000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10100110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10100100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10100000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b10011111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10011110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10011100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10011000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10010111 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10010110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010101 : v_dec_pc_add_3 = (pred_pc + 32'b1110);
	    8'b10010100 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10010000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    8'b10001111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001110 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10001011 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001010 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001001 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10001000 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000111 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10000110 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000101 : v_dec_pc_add_3 = (pred_pc + 32'b1100);
	    8'b10000100 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000011 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000010 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000001 : v_dec_pc_add_3 = (pred_pc + 32'b1010);
	    8'b10000000 : v_dec_pc_add_3 = (pred_pc + 32'b1000);
	    default : v_dec_pc_add_3 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111110 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1111100 : v_dec_inst_4 = data[127:96];
	    8'b1111011 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1111010 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1111001 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1111000 : v_dec_inst_4 = data[111:80];
	    8'b1110110 : v_dec_inst_4 = data[127:96];
	    8'b1110100 : v_dec_inst_4 = data[127:96];
	    8'b1110011 : v_dec_inst_4 = data[127:96];
	    8'b1110010 : v_dec_inst_4 = data[127:96];
	    8'b1110001 : v_dec_inst_4 = data[127:96];
	    8'b1110000 : v_dec_inst_4 = data[95:64];
	    8'b1101111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101110 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101100 : v_dec_inst_4 = data[111:80];
	    8'b1101011 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101010 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101001 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1101000 : v_dec_inst_4 = data[111:80];
	    8'b1100111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1100110 : v_dec_inst_4 = data[111:80];
	    8'b1100101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b1100100 : v_dec_inst_4 = data[111:80];
	    8'b1100011 : v_dec_inst_4 = data[111:80];
	    8'b1100010 : v_dec_inst_4 = data[111:80];
	    8'b1100001 : v_dec_inst_4 = data[111:80];
	    8'b1100000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b1011110 : v_dec_inst_4 = data[127:96];
	    8'b1011100 : v_dec_inst_4 = data[127:96];
	    8'b1011011 : v_dec_inst_4 = data[127:96];
	    8'b1011010 : v_dec_inst_4 = data[127:96];
	    8'b1011001 : v_dec_inst_4 = data[127:96];
	    8'b1011000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1010110 : v_dec_inst_4 = data[127:96];
	    8'b1010100 : v_dec_inst_4 = data[127:96];
	    8'b1010011 : v_dec_inst_4 = data[127:96];
	    8'b1010010 : v_dec_inst_4 = data[127:96];
	    8'b1010001 : v_dec_inst_4 = data[127:96];
	    8'b1010000 : v_dec_inst_4 = data[95:64];
	    8'b1001111 : v_dec_inst_4 = data[127:96];
	    8'b1001110 : v_dec_inst_4 = data[127:96];
	    8'b1001101 : v_dec_inst_4 = data[127:96];
	    8'b1001100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1001011 : v_dec_inst_4 = data[127:96];
	    8'b1001010 : v_dec_inst_4 = data[127:96];
	    8'b1001001 : v_dec_inst_4 = data[127:96];
	    8'b1001000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000111 : v_dec_inst_4 = data[127:96];
	    8'b1000110 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000101 : v_dec_inst_4 = data[127:96];
	    8'b1000100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000011 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000010 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000001 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1000000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b111111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111110 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b111011 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111010 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111001 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b111000 : v_dec_inst_4 = data[111:80];
	    8'b110111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b110110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b110100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110000 : v_dec_inst_4 = data[95:64];
	    8'b101111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101110 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101100 : v_dec_inst_4 = data[111:80];
	    8'b101011 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101010 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101001 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b101000 : v_dec_inst_4 = data[111:80];
	    8'b100111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b100110 : v_dec_inst_4 = data[111:80];
	    8'b100101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b100100 : v_dec_inst_4 = data[111:80];
	    8'b100011 : v_dec_inst_4 = data[111:80];
	    8'b100010 : v_dec_inst_4 = data[111:80];
	    8'b100001 : v_dec_inst_4 = data[111:80];
	    8'b100000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b11111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b11110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b11101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b11100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b11011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b11010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b11001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b11000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10111 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b10110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10101 : v_dec_inst_4 = {16'b0, data[127:112]};
	    8'b10100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10000 : v_dec_inst_4 = data[95:64];
	    8'b1111 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1101 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b1000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b111 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b110 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b101 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b1 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b0 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b11111110 : v_dec_inst_4 = data[143:112];
	    8'b11111100 : v_dec_inst_4 = data[127:96];
	    8'b11111011 : v_dec_inst_4 = data[143:112];
	    8'b11111010 : v_dec_inst_4 = data[143:112];
	    8'b11111001 : v_dec_inst_4 = data[143:112];
	    8'b11111000 : v_dec_inst_4 = data[111:80];
	    8'b11110110 : v_dec_inst_4 = data[127:96];
	    8'b11110100 : v_dec_inst_4 = data[127:96];
	    8'b11110011 : v_dec_inst_4 = data[127:96];
	    8'b11110010 : v_dec_inst_4 = data[127:96];
	    8'b11110001 : v_dec_inst_4 = data[127:96];
	    8'b11110000 : v_dec_inst_4 = data[95:64];
	    8'b11101111 : v_dec_inst_4 = data[143:112];
	    8'b11101110 : v_dec_inst_4 = data[143:112];
	    8'b11101101 : v_dec_inst_4 = data[143:112];
	    8'b11101100 : v_dec_inst_4 = data[111:80];
	    8'b11101011 : v_dec_inst_4 = data[143:112];
	    8'b11101010 : v_dec_inst_4 = data[143:112];
	    8'b11101001 : v_dec_inst_4 = data[143:112];
	    8'b11101000 : v_dec_inst_4 = data[111:80];
	    8'b11100111 : v_dec_inst_4 = data[143:112];
	    8'b11100110 : v_dec_inst_4 = data[111:80];
	    8'b11100101 : v_dec_inst_4 = data[143:112];
	    8'b11100100 : v_dec_inst_4 = data[111:80];
	    8'b11100011 : v_dec_inst_4 = data[111:80];
	    8'b11100010 : v_dec_inst_4 = data[111:80];
	    8'b11100001 : v_dec_inst_4 = data[111:80];
	    8'b11100000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b11011110 : v_dec_inst_4 = data[127:96];
	    8'b11011100 : v_dec_inst_4 = data[127:96];
	    8'b11011011 : v_dec_inst_4 = data[127:96];
	    8'b11011010 : v_dec_inst_4 = data[127:96];
	    8'b11011001 : v_dec_inst_4 = data[127:96];
	    8'b11011000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11010110 : v_dec_inst_4 = data[127:96];
	    8'b11010100 : v_dec_inst_4 = data[127:96];
	    8'b11010011 : v_dec_inst_4 = data[127:96];
	    8'b11010010 : v_dec_inst_4 = data[127:96];
	    8'b11010001 : v_dec_inst_4 = data[127:96];
	    8'b11010000 : v_dec_inst_4 = data[95:64];
	    8'b11001111 : v_dec_inst_4 = data[127:96];
	    8'b11001110 : v_dec_inst_4 = data[127:96];
	    8'b11001101 : v_dec_inst_4 = data[127:96];
	    8'b11001100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11001011 : v_dec_inst_4 = data[127:96];
	    8'b11001010 : v_dec_inst_4 = data[127:96];
	    8'b11001001 : v_dec_inst_4 = data[127:96];
	    8'b11001000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000111 : v_dec_inst_4 = data[127:96];
	    8'b11000110 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000101 : v_dec_inst_4 = data[127:96];
	    8'b11000100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000011 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000010 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000001 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b11000000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b10111111 : v_dec_inst_4 = data[143:112];
	    8'b10111110 : v_dec_inst_4 = data[143:112];
	    8'b10111101 : v_dec_inst_4 = data[143:112];
	    8'b10111100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10111011 : v_dec_inst_4 = data[143:112];
	    8'b10111010 : v_dec_inst_4 = data[143:112];
	    8'b10111001 : v_dec_inst_4 = data[143:112];
	    8'b10111000 : v_dec_inst_4 = data[111:80];
	    8'b10110111 : v_dec_inst_4 = data[143:112];
	    8'b10110110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10110101 : v_dec_inst_4 = data[143:112];
	    8'b10110100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10110011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10110010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10110001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10110000 : v_dec_inst_4 = data[95:64];
	    8'b10101111 : v_dec_inst_4 = data[143:112];
	    8'b10101110 : v_dec_inst_4 = data[143:112];
	    8'b10101101 : v_dec_inst_4 = data[143:112];
	    8'b10101100 : v_dec_inst_4 = data[111:80];
	    8'b10101011 : v_dec_inst_4 = data[143:112];
	    8'b10101010 : v_dec_inst_4 = data[143:112];
	    8'b10101001 : v_dec_inst_4 = data[143:112];
	    8'b10101000 : v_dec_inst_4 = data[111:80];
	    8'b10100111 : v_dec_inst_4 = data[143:112];
	    8'b10100110 : v_dec_inst_4 = data[111:80];
	    8'b10100101 : v_dec_inst_4 = data[143:112];
	    8'b10100100 : v_dec_inst_4 = data[111:80];
	    8'b10100011 : v_dec_inst_4 = data[111:80];
	    8'b10100010 : v_dec_inst_4 = data[111:80];
	    8'b10100001 : v_dec_inst_4 = data[111:80];
	    8'b10100000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    8'b10011111 : v_dec_inst_4 = data[143:112];
	    8'b10011110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011101 : v_dec_inst_4 = data[143:112];
	    8'b10011100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10011000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10010111 : v_dec_inst_4 = data[143:112];
	    8'b10010110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010101 : v_dec_inst_4 = data[143:112];
	    8'b10010100 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10010000 : v_dec_inst_4 = data[95:64];
	    8'b10001111 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001110 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001101 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10001011 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001010 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001001 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10001000 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000111 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10000110 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000101 : v_dec_inst_4 = {16'b0, data[111:96]};
	    8'b10000100 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000011 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000010 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000001 : v_dec_inst_4 = {16'b0, data[95:80]};
	    8'b10000000 : v_dec_inst_4 = {16'b0, data[79:64]};
	    default : v_dec_inst_4 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111110 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1111100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1111011 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1111010 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1111001 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1111000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1110110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1110100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1110011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1110010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1110001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1110000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b1101111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101110 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1101011 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101010 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101001 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1101000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1100110 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b1100100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100011 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100010 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100001 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b1100000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b1011110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1011100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1011011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1011010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1011001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1011000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1010110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1010100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1010011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1010010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1010001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1010000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b1001111 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001101 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1001011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1001000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000111 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1000110 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000101 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b1000100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000011 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000010 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000001 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1000000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b111111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111110 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b111011 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111010 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111001 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b111000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b110111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b110110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b110100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b101111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101110 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b101011 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101010 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101001 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b101000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b100110 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b100100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100011 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100010 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100001 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b100000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b11111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b11110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b11101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b11100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b11011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b11010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b11001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b11000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10111 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b10110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10101 : v_dec_ena_4 = (v_ena[7] && v_vld[7]);
	    8'b10100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b1111 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1101 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b1000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b111 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b110 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b101 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b1 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b0 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b11111110 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11111100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11111011 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11111010 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11111001 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11111000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11110110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11110100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11110011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11110010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11110001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11110000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b11101111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101110 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11101011 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101010 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101001 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11101000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11100110 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b11100100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100011 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100010 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100001 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b11100000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b11011110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11011100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11011011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11011010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11011001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11011000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11010110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11010100 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11010011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11010010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11010001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11010000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b11001111 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001110 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001101 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11001011 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001010 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001001 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11001000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000111 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11000110 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000101 : v_dec_ena_4 = (v_ena[6] && v_vld[7]);
	    8'b11000100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000011 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000010 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000001 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b11000000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b10111111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111110 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10111011 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111010 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111001 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10111000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10110111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10110110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10110101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10110100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10110011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10110010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10110001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10110000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b10101111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101110 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10101011 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101010 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101001 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10101000 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10100110 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10100100 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100011 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100010 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100001 : v_dec_ena_4 = (v_ena[5] && v_vld[6]);
	    8'b10100000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    8'b10011111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10011110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10011100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10011000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10010111 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10010110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010101 : v_dec_ena_4 = (v_ena[7] && v_vld[8]);
	    8'b10010100 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10010000 : v_dec_ena_4 = (v_ena[4] && v_vld[5]);
	    8'b10001111 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001110 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001101 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10001011 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001010 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001001 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10001000 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000111 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10000110 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000101 : v_dec_ena_4 = (v_ena[6] && v_vld[6]);
	    8'b10000100 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000011 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000010 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000001 : v_dec_ena_4 = (v_ena[5] && v_vld[5]);
	    8'b10000000 : v_dec_ena_4 = (v_ena[4] && v_vld[4]);
	    default : v_dec_ena_4 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1111100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1111011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1111010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1111001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1111000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1110110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1110000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1101111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1101011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1100000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b1011110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1011000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1010110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1001111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1001011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1000000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b111111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b111011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b110111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b101111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b101011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b100000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b1111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b1 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b0 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11111110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11111100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11111011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11111010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11111001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11111000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11110110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11110000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11101111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11101011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11100000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b11011110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11011000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11010110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b11001111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11001011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11000000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10111111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10111011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10110111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10101111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101110 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10101011 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101010 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101001 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10100000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    8'b10011111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10011000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10010111 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010101 : v_dec_vld_4 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010100 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[5]));
	    8'b10001111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001110 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10001011 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001010 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001001 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001000 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000111 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000110 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000101 : v_dec_vld_4 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000100 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000011 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000010 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000001 : v_dec_vld_4 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10000000 : v_dec_vld_4 = (v_ena[4] && (v_ena[4] ^ v_vld[4]));
	    default : v_dec_vld_4 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1111100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1111011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1111010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1111001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1111000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1110110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1110100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1110011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1110010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1110001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1110000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1101111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1101011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1101000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1100110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1100100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b1011110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1011100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1011011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1011010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1011001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1011000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1010110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1010100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1010011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1010010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1010001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1010000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1001111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1001011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1001000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1000110 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b1000100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000011 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000010 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000001 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1000000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b111111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b111011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b111000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b110110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b110100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b101111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b101011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b101000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b100110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b100100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b11111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b10110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b10100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1111 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1101 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b1000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b111 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b110 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b101 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b1 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b0 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b11111110 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11111100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11111011 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11111010 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11111001 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11111000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11110110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11110000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11101111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101110 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11101011 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101010 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101001 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11101000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11100110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b11100100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b11100000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b11011110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11011100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11011011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11011010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11011001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11011000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11010110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11010100 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11010011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11010010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11010001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11010000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11001111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001110 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11001011 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001010 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001001 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11001000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000111 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11000110 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000101 : v_dec_pc_add_4 = (pred_pc + 32'b10000);
	    8'b11000100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000011 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000010 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000001 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b11000000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b10111111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111110 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10111011 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111010 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111001 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10111000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10110110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10110100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10110000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10101111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101110 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10101011 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101010 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101001 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10101000 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10100110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10100100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10100000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    8'b10011111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10011110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10011100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10011000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10010111 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10010110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010101 : v_dec_pc_add_4 = (pred_pc + 32'b10010);
	    8'b10010100 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10010000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10001111 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001110 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001101 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10001011 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001010 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001001 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10001000 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000111 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10000110 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000101 : v_dec_pc_add_4 = (pred_pc + 32'b1110);
	    8'b10000100 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000011 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000010 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000001 : v_dec_pc_add_4 = (pred_pc + 32'b1100);
	    8'b10000000 : v_dec_pc_add_4 = (pred_pc + 32'b1010);
	    default : v_dec_pc_add_4 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111000 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1110000 : v_dec_inst_5 = data[127:96];
	    8'b1101100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1101000 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100000 : v_dec_inst_5 = data[111:80];
	    8'b1011000 : v_dec_inst_5 = data[127:96];
	    8'b1010000 : v_dec_inst_5 = data[127:96];
	    8'b1001100 : v_dec_inst_5 = data[127:96];
	    8'b1001000 : v_dec_inst_5 = data[127:96];
	    8'b1000110 : v_dec_inst_5 = data[127:96];
	    8'b1000100 : v_dec_inst_5 = data[127:96];
	    8'b1000011 : v_dec_inst_5 = data[127:96];
	    8'b1000010 : v_dec_inst_5 = data[127:96];
	    8'b1000001 : v_dec_inst_5 = data[127:96];
	    8'b1000000 : v_dec_inst_5 = {16'b0, data[95:80]};
	    8'b111100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b111000 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b101100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b101000 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100000 : v_dec_inst_5 = data[111:80];
	    8'b11110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b11100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b11011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b11010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b11001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b11000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b10100 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b10011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b10010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b10001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b10000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b1111 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1110 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1101 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1100 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b1011 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1010 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1001 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b1000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b111 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b110 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b101 : v_dec_inst_5 = {16'b0, data[127:112]};
	    8'b100 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b11 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b1 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b0 : v_dec_inst_5 = {16'b0, data[95:80]};
	    8'b11111000 : v_dec_inst_5 = data[143:112];
	    8'b11110000 : v_dec_inst_5 = data[127:96];
	    8'b11101100 : v_dec_inst_5 = data[143:112];
	    8'b11101000 : v_dec_inst_5 = data[143:112];
	    8'b11100110 : v_dec_inst_5 = data[143:112];
	    8'b11100100 : v_dec_inst_5 = data[143:112];
	    8'b11100011 : v_dec_inst_5 = data[143:112];
	    8'b11100010 : v_dec_inst_5 = data[143:112];
	    8'b11100001 : v_dec_inst_5 = data[143:112];
	    8'b11100000 : v_dec_inst_5 = data[111:80];
	    8'b11011000 : v_dec_inst_5 = data[127:96];
	    8'b11010000 : v_dec_inst_5 = data[127:96];
	    8'b11001100 : v_dec_inst_5 = data[127:96];
	    8'b11001000 : v_dec_inst_5 = data[127:96];
	    8'b11000110 : v_dec_inst_5 = data[127:96];
	    8'b11000100 : v_dec_inst_5 = data[127:96];
	    8'b11000011 : v_dec_inst_5 = data[127:96];
	    8'b11000010 : v_dec_inst_5 = data[127:96];
	    8'b11000001 : v_dec_inst_5 = data[127:96];
	    8'b11000000 : v_dec_inst_5 = {16'b0, data[95:80]};
	    8'b10111100 : v_dec_inst_5 = data[143:112];
	    8'b10111000 : v_dec_inst_5 = data[143:112];
	    8'b10110110 : v_dec_inst_5 = data[143:112];
	    8'b10110100 : v_dec_inst_5 = data[143:112];
	    8'b10110011 : v_dec_inst_5 = data[143:112];
	    8'b10110010 : v_dec_inst_5 = data[143:112];
	    8'b10110001 : v_dec_inst_5 = data[143:112];
	    8'b10110000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10101100 : v_dec_inst_5 = data[143:112];
	    8'b10101000 : v_dec_inst_5 = data[143:112];
	    8'b10100110 : v_dec_inst_5 = data[143:112];
	    8'b10100100 : v_dec_inst_5 = data[143:112];
	    8'b10100011 : v_dec_inst_5 = data[143:112];
	    8'b10100010 : v_dec_inst_5 = data[143:112];
	    8'b10100001 : v_dec_inst_5 = data[143:112];
	    8'b10100000 : v_dec_inst_5 = data[111:80];
	    8'b10011110 : v_dec_inst_5 = data[143:112];
	    8'b10011100 : v_dec_inst_5 = data[143:112];
	    8'b10011011 : v_dec_inst_5 = data[143:112];
	    8'b10011010 : v_dec_inst_5 = data[143:112];
	    8'b10011001 : v_dec_inst_5 = data[143:112];
	    8'b10011000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10010110 : v_dec_inst_5 = data[143:112];
	    8'b10010100 : v_dec_inst_5 = data[143:112];
	    8'b10010011 : v_dec_inst_5 = data[143:112];
	    8'b10010010 : v_dec_inst_5 = data[143:112];
	    8'b10010001 : v_dec_inst_5 = data[143:112];
	    8'b10010000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10001111 : v_dec_inst_5 = data[143:112];
	    8'b10001110 : v_dec_inst_5 = data[143:112];
	    8'b10001101 : v_dec_inst_5 = data[143:112];
	    8'b10001100 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10001011 : v_dec_inst_5 = data[143:112];
	    8'b10001010 : v_dec_inst_5 = data[143:112];
	    8'b10001001 : v_dec_inst_5 = data[143:112];
	    8'b10001000 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000111 : v_dec_inst_5 = data[143:112];
	    8'b10000110 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000101 : v_dec_inst_5 = data[143:112];
	    8'b10000100 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000011 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000010 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000001 : v_dec_inst_5 = {16'b0, data[111:96]};
	    8'b10000000 : v_dec_inst_5 = {16'b0, data[95:80]};
	    default : v_dec_inst_5 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111000 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1110000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1101100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1101000 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100000 : v_dec_ena_5 = (v_ena[5] && v_vld[6]);
	    8'b1011000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1010000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1001100 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1001000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000110 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000100 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000011 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000010 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000001 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b1000000 : v_dec_ena_5 = (v_ena[5] && v_vld[5]);
	    8'b111100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b111000 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b101100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b101000 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100000 : v_dec_ena_5 = (v_ena[5] && v_vld[6]);
	    8'b11110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b11100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b11011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b11010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b11001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b11000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b10100 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b10011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b10010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b10001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b10000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b1111 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1110 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1101 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1100 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b1011 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1010 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1001 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b1000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b111 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b110 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b101 : v_dec_ena_5 = (v_ena[7] && v_vld[7]);
	    8'b100 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b11 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b1 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b0 : v_dec_ena_5 = (v_ena[5] && v_vld[5]);
	    8'b11111000 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11110000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11101100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11101000 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b11100000 : v_dec_ena_5 = (v_ena[5] && v_vld[6]);
	    8'b11011000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11010000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11001100 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11001000 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000110 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000100 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000011 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000010 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000001 : v_dec_ena_5 = (v_ena[6] && v_vld[7]);
	    8'b11000000 : v_dec_ena_5 = (v_ena[5] && v_vld[5]);
	    8'b10111100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10111000 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10110000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10101100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10101000 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10100000 : v_dec_ena_5 = (v_ena[5] && v_vld[6]);
	    8'b10011110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10011100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10011011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10011010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10011001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10011000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10010110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10010100 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10010011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10010010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10010001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10010000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10001111 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001110 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001101 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001100 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10001011 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001010 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001001 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10001000 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000111 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10000110 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000101 : v_dec_ena_5 = (v_ena[7] && v_vld[8]);
	    8'b10000100 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000011 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000010 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000001 : v_dec_ena_5 = (v_ena[6] && v_vld[6]);
	    8'b10000000 : v_dec_ena_5 = (v_ena[5] && v_vld[5]);
	    default : v_dec_ena_5 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1110000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1101100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b1011000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1010000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1001000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000110 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000011 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000010 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000001 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b1000000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b111100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b111000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b101100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b101000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1111 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1101 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b111 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b101 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b1 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b0 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b11111000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11110000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11101100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11101000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11100000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b11011000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11010000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11001000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000110 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000011 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000010 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000001 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b11000000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    8'b10111100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10111000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10110000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10101100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10101000 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[6]));
	    8'b10011110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10010110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010100 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001111 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001110 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001101 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10001011 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001010 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001001 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001000 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000111 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000110 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000101 : v_dec_vld_5 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000100 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000011 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000010 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000001 : v_dec_vld_5 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b10000000 : v_dec_vld_5 = (v_ena[5] && (v_ena[5] ^ v_vld[5]));
	    default : v_dec_vld_5 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1111000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1110000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1101100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1101000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b1011000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1010000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1001100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1001000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000000 : v_dec_pc_add_5 = (pred_pc + 32'b1100);
	    8'b111100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b111000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b101100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b101000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b11110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b10100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b10011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b10010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b10001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b10000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b1111 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1101 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1100 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b1011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b1000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b111 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b110 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b101 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b100 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b11 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b1 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b0 : v_dec_pc_add_5 = (pred_pc + 32'b1100);
	    8'b11111000 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11110000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11101100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11101000 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b11100000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b11011000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11010000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11001100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11001000 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000110 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000100 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000011 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000010 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000001 : v_dec_pc_add_5 = (pred_pc + 32'b10000);
	    8'b11000000 : v_dec_pc_add_5 = (pred_pc + 32'b1100);
	    8'b10111100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10111000 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10110000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10101100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10101000 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10100000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10011110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10011100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10011011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10011010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10011001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10011000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10010110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10010100 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10010011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10010010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10010001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10010000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10001111 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001110 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001101 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001100 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10001011 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001010 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001001 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10001000 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000111 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10000110 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000101 : v_dec_pc_add_5 = (pred_pc + 32'b10010);
	    8'b10000100 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000011 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000010 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000001 : v_dec_pc_add_5 = (pred_pc + 32'b1110);
	    8'b10000000 : v_dec_pc_add_5 = (pred_pc + 32'b1100);
	    default : v_dec_pc_add_5 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1100000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b1000000 : v_dec_inst_6 = data[127:96];
	    8'b110000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b100000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b11000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b10000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b1100 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b1000 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b110 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b100 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b11 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b10 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b1 : v_dec_inst_6 = {16'b0, data[127:112]};
	    8'b0 : v_dec_inst_6 = {16'b0, data[111:96]};
	    8'b11100000 : v_dec_inst_6 = data[143:112];
	    8'b11000000 : v_dec_inst_6 = data[127:96];
	    8'b10110000 : v_dec_inst_6 = data[143:112];
	    8'b10100000 : v_dec_inst_6 = data[143:112];
	    8'b10011000 : v_dec_inst_6 = data[143:112];
	    8'b10010000 : v_dec_inst_6 = data[143:112];
	    8'b10001100 : v_dec_inst_6 = data[143:112];
	    8'b10001000 : v_dec_inst_6 = data[143:112];
	    8'b10000110 : v_dec_inst_6 = data[143:112];
	    8'b10000100 : v_dec_inst_6 = data[143:112];
	    8'b10000011 : v_dec_inst_6 = data[143:112];
	    8'b10000010 : v_dec_inst_6 = data[143:112];
	    8'b10000001 : v_dec_inst_6 = data[143:112];
	    8'b10000000 : v_dec_inst_6 = {16'b0, data[111:96]};
	    default : v_dec_inst_6 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1100000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b1000000 : v_dec_ena_6 = (v_ena[6] && v_vld[7]);
	    8'b110000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b100000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b11000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b10000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b1100 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b1000 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b110 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b100 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b11 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b10 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b1 : v_dec_ena_6 = (v_ena[7] && v_vld[7]);
	    8'b0 : v_dec_ena_6 = (v_ena[6] && v_vld[6]);
	    8'b11100000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b11000000 : v_dec_ena_6 = (v_ena[6] && v_vld[7]);
	    8'b10110000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10100000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10011000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10010000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10001100 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10001000 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000110 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000100 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000011 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000010 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000001 : v_dec_ena_6 = (v_ena[7] && v_vld[8]);
	    8'b10000000 : v_dec_ena_6 = (v_ena[6] && v_vld[6]);
	    default : v_dec_ena_6 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1100000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1000000 : v_dec_vld_6 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b110000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1100 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b110 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b100 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b11 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b1 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b0 : v_dec_vld_6 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    8'b11100000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b11000000 : v_dec_vld_6 = (v_ena[6] && (v_ena[6] ^ v_vld[7]));
	    8'b10110000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10100000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10011000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10010000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001100 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10001000 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000110 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000100 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000011 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000010 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000001 : v_dec_vld_6 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    8'b10000000 : v_dec_vld_6 = (v_ena[6] && (v_ena[6] ^ v_vld[6]));
	    default : v_dec_vld_6 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b1100000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b1000000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b110000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b100000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b11000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b10000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b1100 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b1000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b110 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b100 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b11 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b10 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b1 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b0 : v_dec_pc_add_6 = (pred_pc + 32'b1110);
	    8'b11100000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b11000000 : v_dec_pc_add_6 = (pred_pc + 32'b10000);
	    8'b10110000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10100000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10011000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10010000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10001100 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10001000 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000110 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000100 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000011 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000010 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000001 : v_dec_pc_add_6 = (pred_pc + 32'b10010);
	    8'b10000000 : v_dec_pc_add_6 = (pred_pc + 32'b1110);
	    default : v_dec_pc_add_6 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b0 : v_dec_inst_7 = {16'b0, data[127:112]};
	    8'b10000000 : v_dec_inst_7 = data[143:112];
	    default : v_dec_inst_7 = 32'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b0 : v_dec_ena_7 = (v_ena[7] && v_vld[7]);
	    8'b10000000 : v_dec_ena_7 = (v_ena[7] && v_vld[8]);
	    default : v_dec_ena_7 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b0 : v_dec_vld_7 = (v_ena[7] && (v_ena[7] ^ v_vld[7]));
	    8'b10000000 : v_dec_vld_7 = (v_ena[7] && (v_ena[7] ^ v_vld[8]));
	    default : v_dec_vld_7 = 1'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b0 : v_dec_pc_add_7 = (pred_pc + 32'b10000);
	    8'b10000000 : v_dec_pc_add_7 = (pred_pc + 32'b10010);
	    default : v_dec_pc_add_7 = 33'b0;
	    endcase
	end
	
	always @(*) begin
	    case(v_inst_type[7:0])
	    8'b11111110 : use_last_w = 1'b1;
	    8'b11111011 : use_last_w = 1'b1;
	    8'b11111010 : use_last_w = 1'b1;
	    8'b11111001 : use_last_w = 1'b1;
	    8'b11101111 : use_last_w = 1'b1;
	    8'b11101110 : use_last_w = 1'b1;
	    8'b11101101 : use_last_w = 1'b1;
	    8'b11101011 : use_last_w = 1'b1;
	    8'b11101010 : use_last_w = 1'b1;
	    8'b11101001 : use_last_w = 1'b1;
	    8'b11100111 : use_last_w = 1'b1;
	    8'b11100101 : use_last_w = 1'b1;
	    8'b10111111 : use_last_w = 1'b1;
	    8'b10111110 : use_last_w = 1'b1;
	    8'b10111101 : use_last_w = 1'b1;
	    8'b10111011 : use_last_w = 1'b1;
	    8'b10111010 : use_last_w = 1'b1;
	    8'b10111001 : use_last_w = 1'b1;
	    8'b10110111 : use_last_w = 1'b1;
	    8'b10110101 : use_last_w = 1'b1;
	    8'b10101111 : use_last_w = 1'b1;
	    8'b10101110 : use_last_w = 1'b1;
	    8'b10101101 : use_last_w = 1'b1;
	    8'b10101011 : use_last_w = 1'b1;
	    8'b10101010 : use_last_w = 1'b1;
	    8'b10101001 : use_last_w = 1'b1;
	    8'b10100111 : use_last_w = 1'b1;
	    8'b10100101 : use_last_w = 1'b1;
	    8'b10011111 : use_last_w = 1'b1;
	    8'b10011101 : use_last_w = 1'b1;
	    8'b10010111 : use_last_w = 1'b1;
	    8'b10010101 : use_last_w = 1'b1;
	    8'b11111000 : use_last_w = 1'b1;
	    8'b11101100 : use_last_w = 1'b1;
	    8'b11101000 : use_last_w = 1'b1;
	    8'b11100110 : use_last_w = 1'b1;
	    8'b11100100 : use_last_w = 1'b1;
	    8'b11100011 : use_last_w = 1'b1;
	    8'b11100010 : use_last_w = 1'b1;
	    8'b11100001 : use_last_w = 1'b1;
	    8'b10111100 : use_last_w = 1'b1;
	    8'b10111000 : use_last_w = 1'b1;
	    8'b10110110 : use_last_w = 1'b1;
	    8'b10110100 : use_last_w = 1'b1;
	    8'b10110011 : use_last_w = 1'b1;
	    8'b10110010 : use_last_w = 1'b1;
	    8'b10110001 : use_last_w = 1'b1;
	    8'b10101100 : use_last_w = 1'b1;
	    8'b10101000 : use_last_w = 1'b1;
	    8'b10100110 : use_last_w = 1'b1;
	    8'b10100100 : use_last_w = 1'b1;
	    8'b10100011 : use_last_w = 1'b1;
	    8'b10100010 : use_last_w = 1'b1;
	    8'b10100001 : use_last_w = 1'b1;
	    8'b10011110 : use_last_w = 1'b1;
	    8'b10011100 : use_last_w = 1'b1;
	    8'b10011011 : use_last_w = 1'b1;
	    8'b10011010 : use_last_w = 1'b1;
	    8'b10011001 : use_last_w = 1'b1;
	    8'b10010110 : use_last_w = 1'b1;
	    8'b10010100 : use_last_w = 1'b1;
	    8'b10010011 : use_last_w = 1'b1;
	    8'b10010010 : use_last_w = 1'b1;
	    8'b10010001 : use_last_w = 1'b1;
	    8'b10001111 : use_last_w = 1'b1;
	    8'b10001110 : use_last_w = 1'b1;
	    8'b10001101 : use_last_w = 1'b1;
	    8'b10001011 : use_last_w = 1'b1;
	    8'b10001010 : use_last_w = 1'b1;
	    8'b10001001 : use_last_w = 1'b1;
	    8'b10000111 : use_last_w = 1'b1;
	    8'b10000101 : use_last_w = 1'b1;
	    8'b11100000 : use_last_w = 1'b1;
	    8'b10110000 : use_last_w = 1'b1;
	    8'b10100000 : use_last_w = 1'b1;
	    8'b10011000 : use_last_w = 1'b1;
	    8'b10010000 : use_last_w = 1'b1;
	    8'b10001100 : use_last_w = 1'b1;
	    8'b10001000 : use_last_w = 1'b1;
	    8'b10000110 : use_last_w = 1'b1;
	    8'b10000100 : use_last_w = 1'b1;
	    8'b10000011 : use_last_w = 1'b1;
	    8'b10000010 : use_last_w = 1'b1;
	    8'b10000001 : use_last_w = 1'b1;
	    8'b10000000 : use_last_w = 1'b1;
	    default : use_last_w = 1'b0;
	    endcase
	end
	

	//Wire this module connect to sub module.

	//module inst.
	cmn_lead_one_rev #(
		.ENTRY_NUM(32'd8))
	u_dec_oh (
		.v_entry_vld(v_dec_ena),
		.v_free_idx_oh(v_dec_last),
		.v_free_idx_bin(),
		.v_free_vld());

endmodule
//[UHDL]Content End [md5:3634c664f0cae32a29033e3a1552312c]

